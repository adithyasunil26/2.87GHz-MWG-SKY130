magic
tech sky130A
timestamp 1647788355
<< psubdiff >>
rect 4315 75 4445 90
rect 4315 -25 4330 75
rect 4430 -25 4445 75
rect 4315 -40 4445 -25
rect -329 -121 -199 -106
rect -329 -221 -314 -121
rect -214 -221 -199 -121
rect -329 -236 -199 -221
rect 4518 -145 4648 -130
rect 4315 -255 4445 -240
rect 4315 -355 4330 -255
rect 4430 -355 4445 -255
rect 4518 -245 4533 -145
rect 4633 -245 4648 -145
rect 4518 -260 4648 -245
rect 4315 -370 4445 -355
rect 4315 -585 4445 -570
rect -329 -611 -199 -596
rect -329 -711 -314 -611
rect -214 -711 -199 -611
rect 4315 -685 4330 -585
rect 4430 -685 4445 -585
rect 4315 -700 4445 -685
rect 4518 -635 4648 -620
rect -329 -726 -199 -711
rect 4518 -735 4533 -635
rect 4633 -735 4648 -635
rect 4518 -750 4648 -735
rect 4315 -915 4445 -900
rect 4315 -1015 4330 -915
rect 4430 -1015 4445 -915
rect 4315 -1030 4445 -1015
rect -329 -1101 -199 -1086
rect -329 -1201 -314 -1101
rect -214 -1201 -199 -1101
rect -329 -1216 -199 -1201
rect 4518 -1125 4648 -1110
rect 4518 -1225 4533 -1125
rect 4633 -1225 4648 -1125
rect 4315 -1245 4445 -1230
rect 4518 -1240 4648 -1225
rect 4315 -1345 4330 -1245
rect 4430 -1345 4445 -1245
rect 4315 -1360 4445 -1345
rect -329 -1458 -199 -1443
rect -329 -1558 -314 -1458
rect -214 -1558 -199 -1458
rect -329 -1573 -199 -1558
rect 4518 -1482 4648 -1467
rect 4315 -1575 4445 -1560
rect 4315 -1675 4330 -1575
rect 4430 -1675 4445 -1575
rect 4518 -1582 4533 -1482
rect 4633 -1582 4648 -1482
rect 4518 -1597 4648 -1582
rect 4315 -1690 4445 -1675
rect 4315 -1905 4445 -1890
rect -329 -1948 -199 -1933
rect -329 -2048 -314 -1948
rect -214 -2048 -199 -1948
rect 4315 -2005 4330 -1905
rect 4430 -2005 4445 -1905
rect 4315 -2020 4445 -2005
rect 4518 -1972 4648 -1957
rect -329 -2063 -199 -2048
rect 4518 -2072 4533 -1972
rect 4633 -2072 4648 -1972
rect 4518 -2087 4648 -2072
rect 4315 -2235 4445 -2220
rect 4315 -2335 4330 -2235
rect 4430 -2335 4445 -2235
rect 4315 -2350 4445 -2335
rect -329 -2438 -199 -2423
rect -329 -2538 -314 -2438
rect -214 -2538 -199 -2438
rect -329 -2553 -199 -2538
rect 4518 -2462 4648 -2447
rect 4315 -2565 4445 -2550
rect 4315 -2665 4330 -2565
rect 4430 -2665 4445 -2565
rect 4518 -2562 4533 -2462
rect 4633 -2562 4648 -2462
rect 4518 -2577 4648 -2562
rect 4315 -2680 4445 -2665
rect -329 -2803 -199 -2788
rect -329 -2903 -314 -2803
rect -214 -2903 -199 -2803
rect 4518 -2827 4648 -2812
rect -329 -2918 -199 -2903
rect 4315 -2895 4445 -2880
rect 4315 -2995 4330 -2895
rect 4430 -2995 4445 -2895
rect 4518 -2927 4533 -2827
rect 4633 -2927 4648 -2827
rect 4518 -2942 4648 -2927
rect 4315 -3010 4445 -2995
rect 4315 -3225 4445 -3210
rect -329 -3293 -199 -3278
rect -329 -3393 -314 -3293
rect -214 -3393 -199 -3293
rect 4315 -3325 4330 -3225
rect 4430 -3325 4445 -3225
rect 4315 -3340 4445 -3325
rect 4518 -3317 4648 -3302
rect -329 -3408 -199 -3393
rect 4518 -3417 4533 -3317
rect 4633 -3417 4648 -3317
rect 4518 -3432 4648 -3417
rect 4315 -3555 4445 -3540
rect 4315 -3655 4330 -3555
rect 4430 -3655 4445 -3555
rect 4315 -3670 4445 -3655
rect -329 -3783 -199 -3768
rect -329 -3883 -314 -3783
rect -214 -3883 -199 -3783
rect 4518 -3807 4648 -3792
rect -329 -3898 -199 -3883
rect 4315 -3885 4445 -3870
rect 4315 -3985 4330 -3885
rect 4430 -3985 4445 -3885
rect 4518 -3907 4533 -3807
rect 4633 -3907 4648 -3807
rect 4518 -3922 4648 -3907
rect 4315 -4000 4445 -3985
rect -329 -4148 -199 -4133
rect -329 -4248 -314 -4148
rect -214 -4248 -199 -4148
rect 4518 -4172 4648 -4157
rect -329 -4263 -199 -4248
rect 4315 -4215 4445 -4200
rect 4315 -4315 4330 -4215
rect 4430 -4315 4445 -4215
rect 4518 -4272 4533 -4172
rect 4633 -4272 4648 -4172
rect 4518 -4287 4648 -4272
rect 4315 -4330 4445 -4315
rect 4315 -4545 4445 -4530
rect -329 -4638 -199 -4623
rect -329 -4738 -314 -4638
rect -214 -4738 -199 -4638
rect 4315 -4645 4330 -4545
rect 4430 -4645 4445 -4545
rect 4315 -4660 4445 -4645
rect -329 -4753 -199 -4738
rect 4518 -4662 4648 -4647
rect 4518 -4762 4533 -4662
rect 4633 -4762 4648 -4662
rect 4518 -4777 4648 -4762
rect 4315 -4875 4445 -4860
rect 4315 -4975 4330 -4875
rect 4430 -4975 4445 -4875
rect 4315 -4990 4445 -4975
rect -329 -5128 -199 -5113
rect -329 -5228 -314 -5128
rect -214 -5228 -199 -5128
rect 4518 -5152 4648 -5137
rect -329 -5243 -199 -5228
rect 3895 -5205 4025 -5190
rect 3895 -5305 3910 -5205
rect 4010 -5305 4025 -5205
rect 3895 -5320 4025 -5305
rect 4315 -5205 4445 -5190
rect 4315 -5305 4330 -5205
rect 4430 -5305 4445 -5205
rect 4518 -5252 4533 -5152
rect 4633 -5252 4648 -5152
rect 4518 -5267 4648 -5252
rect 4315 -5320 4445 -5305
rect -204 -5562 -74 -5547
rect -204 -5662 -189 -5562
rect -89 -5662 -74 -5562
rect -204 -5677 -74 -5662
rect 286 -5562 416 -5547
rect 286 -5662 301 -5562
rect 401 -5662 416 -5562
rect 286 -5677 416 -5662
rect 4221 -5561 4351 -5546
rect 4221 -5661 4236 -5561
rect 4336 -5661 4351 -5561
rect 4221 -5676 4351 -5661
<< psubdiffcont >>
rect 4330 -25 4430 75
rect -314 -221 -214 -121
rect 4330 -355 4430 -255
rect 4533 -245 4633 -145
rect -314 -711 -214 -611
rect 4330 -685 4430 -585
rect 4533 -735 4633 -635
rect 4330 -1015 4430 -915
rect -314 -1201 -214 -1101
rect 4533 -1225 4633 -1125
rect 4330 -1345 4430 -1245
rect -314 -1558 -214 -1458
rect 4330 -1675 4430 -1575
rect 4533 -1582 4633 -1482
rect -314 -2048 -214 -1948
rect 4330 -2005 4430 -1905
rect 4533 -2072 4633 -1972
rect 4330 -2335 4430 -2235
rect -314 -2538 -214 -2438
rect 4330 -2665 4430 -2565
rect 4533 -2562 4633 -2462
rect -314 -2903 -214 -2803
rect 4330 -2995 4430 -2895
rect 4533 -2927 4633 -2827
rect -314 -3393 -214 -3293
rect 4330 -3325 4430 -3225
rect 4533 -3417 4633 -3317
rect 4330 -3655 4430 -3555
rect -314 -3883 -214 -3783
rect 4330 -3985 4430 -3885
rect 4533 -3907 4633 -3807
rect -314 -4248 -214 -4148
rect 4330 -4315 4430 -4215
rect 4533 -4272 4633 -4172
rect -314 -4738 -214 -4638
rect 4330 -4645 4430 -4545
rect 4533 -4762 4633 -4662
rect 4330 -4975 4430 -4875
rect -314 -5228 -214 -5128
rect 3910 -5305 4010 -5205
rect 4330 -5305 4430 -5205
rect 4533 -5252 4633 -5152
rect -189 -5662 -89 -5562
rect 301 -5662 401 -5562
rect 4236 -5661 4336 -5561
<< locali >>
rect 3720 750 3810 760
rect 665 740 735 750
rect 665 730 675 740
rect 505 700 675 730
rect 665 690 675 700
rect 725 690 735 740
rect 2210 735 2280 745
rect 2210 725 2220 735
rect 2040 695 2220 725
rect 665 680 735 690
rect 2210 685 2220 695
rect 2270 685 2280 735
rect 3720 730 3730 750
rect 3570 700 3730 730
rect 2210 675 2280 685
rect 3720 680 3730 700
rect 3800 680 3810 750
rect 3720 670 3810 680
rect 3595 565 3735 635
rect 3675 535 3735 565
rect 3675 485 3680 535
rect 3730 485 3735 535
rect 3675 480 3735 485
rect 3598 415 3628 426
rect 3598 338 3606 415
rect 3623 338 3628 415
rect 3598 330 3628 338
rect -346 81 295 245
rect 4108 91 4267 132
rect -346 -121 -186 81
rect 4108 75 4661 91
rect 4108 -25 4330 75
rect 4430 -25 4661 75
rect 4108 -42 4661 -25
rect -346 -221 -314 -121
rect -214 -221 -186 -121
rect -346 -611 -186 -221
rect 4501 -145 4661 -42
rect 4501 -245 4533 -145
rect 4633 -245 4661 -145
rect 4320 -255 4440 -245
rect 4320 -355 4330 -255
rect 4430 -355 4440 -255
rect 4320 -365 4440 -355
rect -346 -711 -314 -611
rect -214 -711 -186 -611
rect 4320 -585 4440 -575
rect 4320 -685 4330 -585
rect 4430 -685 4440 -585
rect 4320 -695 4440 -685
rect 4501 -635 4661 -245
rect -346 -1101 -186 -711
rect 4501 -735 4533 -635
rect 4633 -735 4661 -635
rect 958 -840 1143 -805
rect 1462 -840 1632 -805
rect 1936 -840 2121 -805
rect 2426 -840 2606 -805
rect 2917 -840 3097 -805
rect 3428 -840 3693 -805
rect -346 -1201 -314 -1101
rect -214 -1201 -186 -1101
rect -346 -1458 -186 -1201
rect -346 -1558 -314 -1458
rect -214 -1558 -186 -1458
rect -346 -1634 -186 -1558
rect -346 -1764 565 -1634
rect -346 -1948 -186 -1764
rect -346 -2048 -314 -1948
rect -214 -2048 -186 -1948
rect -346 -2438 -186 -2048
rect -346 -2538 -314 -2438
rect -214 -2538 -186 -2438
rect -346 -2803 -186 -2538
rect 1108 -2575 1143 -840
rect 1597 -2575 1632 -840
rect 2086 -2575 2121 -840
rect 2571 -2575 2606 -840
rect 3062 -2575 3097 -840
rect 3658 -2575 3693 -840
rect 4320 -915 4440 -905
rect 4320 -1015 4330 -915
rect 4430 -1015 4440 -915
rect 4320 -1025 4440 -1015
rect 4501 -1125 4661 -735
rect 4501 -1225 4533 -1125
rect 4633 -1225 4661 -1125
rect 4320 -1245 4440 -1235
rect 4320 -1345 4330 -1245
rect 4430 -1345 4440 -1245
rect 4320 -1355 4440 -1345
rect 4501 -1482 4661 -1225
rect 4320 -1575 4440 -1565
rect 4320 -1675 4330 -1575
rect 4430 -1675 4440 -1575
rect 4320 -1685 4440 -1675
rect 4501 -1582 4533 -1482
rect 4633 -1582 4661 -1482
rect 4320 -1905 4440 -1895
rect 4320 -2005 4330 -1905
rect 4430 -2005 4440 -1905
rect 4320 -2015 4440 -2005
rect 4501 -1972 4661 -1582
rect 4501 -2072 4533 -1972
rect 4633 -2072 4661 -1972
rect 4320 -2235 4440 -2225
rect 4320 -2335 4330 -2235
rect 4430 -2335 4440 -2235
rect 4320 -2345 4440 -2335
rect 4501 -2462 4661 -2072
rect 958 -2610 1143 -2575
rect 1462 -2610 1632 -2575
rect 1936 -2610 2121 -2575
rect 2426 -2610 2606 -2575
rect 2917 -2610 3097 -2575
rect 3428 -2610 3693 -2575
rect -346 -2903 -314 -2803
rect -214 -2903 -186 -2803
rect -346 -3293 -186 -2903
rect -346 -3393 -314 -3293
rect -214 -3393 -186 -3293
rect -346 -3404 -186 -3393
rect -346 -3534 563 -3404
rect -346 -3783 -186 -3534
rect -346 -3883 -314 -3783
rect -214 -3883 -186 -3783
rect -346 -4148 -186 -3883
rect -346 -4248 -314 -4148
rect -214 -4248 -186 -4148
rect -346 -4638 -186 -4248
rect 1108 -4360 1143 -2610
rect 1597 -4360 1632 -2610
rect 2086 -4360 2121 -2610
rect 2571 -4360 2606 -2610
rect 3062 -4360 3097 -2610
rect 3658 -4360 3693 -2610
rect 4320 -2565 4440 -2555
rect 4320 -2665 4330 -2565
rect 4430 -2665 4440 -2565
rect 4320 -2675 4440 -2665
rect 4501 -2562 4533 -2462
rect 4633 -2562 4661 -2462
rect 4501 -2827 4661 -2562
rect 4320 -2895 4440 -2885
rect 4320 -2995 4330 -2895
rect 4430 -2995 4440 -2895
rect 4320 -3005 4440 -2995
rect 4501 -2927 4533 -2827
rect 4633 -2927 4661 -2827
rect 4320 -3225 4440 -3215
rect 4320 -3325 4330 -3225
rect 4430 -3325 4440 -3225
rect 4320 -3335 4440 -3325
rect 4501 -3317 4661 -2927
rect 4501 -3417 4533 -3317
rect 4633 -3417 4661 -3317
rect 4320 -3555 4440 -3545
rect 4320 -3655 4330 -3555
rect 4430 -3655 4440 -3555
rect 4320 -3665 4440 -3655
rect 4501 -3807 4661 -3417
rect 4320 -3885 4440 -3875
rect 4320 -3985 4330 -3885
rect 4430 -3985 4440 -3885
rect 4320 -3995 4440 -3985
rect 4501 -3907 4533 -3807
rect 4633 -3907 4661 -3807
rect 4501 -4172 4661 -3907
rect 4320 -4215 4440 -4205
rect 4320 -4315 4330 -4215
rect 4430 -4315 4440 -4215
rect 4320 -4325 4440 -4315
rect 4501 -4272 4533 -4172
rect 4633 -4272 4661 -4172
rect 958 -4395 1143 -4360
rect 1462 -4395 1632 -4360
rect 1936 -4395 2121 -4360
rect 2426 -4395 2606 -4360
rect 2917 -4395 3097 -4360
rect 3428 -4395 3693 -4360
rect -346 -4738 -314 -4638
rect -214 -4738 -186 -4638
rect 4320 -4545 4440 -4535
rect 4320 -4645 4330 -4545
rect 4430 -4645 4440 -4545
rect 4320 -4655 4440 -4645
rect -346 -5128 -186 -4738
rect 4501 -4662 4661 -4272
rect 4501 -4762 4533 -4662
rect 4633 -4762 4661 -4662
rect 4320 -4875 4440 -4865
rect 4320 -4975 4330 -4875
rect 4430 -4975 4440 -4875
rect 4320 -4985 4440 -4975
rect -346 -5228 -314 -5128
rect -214 -5191 -186 -5128
rect 4501 -5152 4661 -4762
rect -214 -5228 567 -5191
rect -346 -5318 567 -5228
rect 3900 -5205 4020 -5195
rect 3900 -5305 3910 -5205
rect 4010 -5305 4020 -5205
rect 3900 -5315 4020 -5305
rect 4320 -5205 4440 -5195
rect 4320 -5305 4330 -5205
rect 4430 -5305 4440 -5205
rect 4320 -5315 4440 -5305
rect 4501 -5252 4533 -5152
rect 4633 -5252 4661 -5152
rect -348 -5321 567 -5318
rect -348 -5530 -185 -5321
rect 4501 -5389 4661 -5252
rect 4501 -5410 4659 -5389
rect 4502 -5529 4659 -5410
rect -348 -5562 731 -5530
rect -348 -5662 -189 -5562
rect -89 -5662 301 -5562
rect 401 -5662 731 -5562
rect -348 -5688 731 -5662
rect 4207 -5561 4659 -5529
rect 4207 -5661 4236 -5561
rect 4336 -5661 4659 -5561
rect 4207 -5687 4659 -5661
rect -348 -5690 -185 -5688
<< viali >>
rect 675 690 725 740
rect 2220 685 2270 735
rect 3730 680 3800 750
rect 3680 485 3730 535
rect 3606 338 3623 415
rect 4330 -25 4430 75
rect 4330 -355 4430 -255
rect 4330 -685 4430 -585
rect 4330 -1015 4430 -915
rect 4330 -1345 4430 -1245
rect 4330 -1675 4430 -1575
rect 4330 -2005 4430 -1905
rect 4330 -2335 4430 -2235
rect 4330 -2665 4430 -2565
rect 4330 -2995 4430 -2895
rect 4330 -3325 4430 -3225
rect 4330 -3655 4430 -3555
rect 4330 -3985 4430 -3885
rect 4330 -4315 4430 -4215
rect 4330 -4645 4430 -4545
rect 4330 -4975 4430 -4875
rect 3910 -5305 4010 -5205
rect 4330 -5305 4430 -5205
<< metal1 >>
rect 3720 750 3810 760
rect 665 740 735 750
rect 665 690 675 740
rect 725 690 735 740
rect 665 680 735 690
rect 2210 735 2280 745
rect 2210 685 2220 735
rect 2270 685 2280 735
rect 2210 675 2280 685
rect 3720 680 3730 750
rect 3800 680 3810 750
rect 3720 670 3810 680
rect 4325 560 4435 565
rect 4325 555 4330 560
rect 3655 535 4330 555
rect 3655 485 3680 535
rect 3730 485 4330 535
rect 3655 465 4330 485
rect 4325 460 4330 465
rect 4430 460 4435 560
rect 4325 455 4435 460
rect 3598 415 3628 426
rect 3598 338 3606 415
rect 3623 338 3628 415
rect 3598 330 3628 338
rect 4320 75 4440 85
rect 4320 -25 4330 75
rect 4430 -25 4440 75
rect 4320 -35 4440 -25
rect 4320 -255 4440 -245
rect 4320 -355 4330 -255
rect 4430 -355 4440 -255
rect 4320 -365 4440 -355
rect 4320 -585 4440 -575
rect 4320 -685 4330 -585
rect 4430 -685 4440 -585
rect 4320 -695 4440 -685
rect 4320 -915 4440 -905
rect 4320 -1015 4330 -915
rect 4430 -1015 4440 -915
rect 4320 -1025 4440 -1015
rect 4320 -1245 4440 -1235
rect 4320 -1345 4330 -1245
rect 4430 -1345 4440 -1245
rect 4320 -1355 4440 -1345
rect 4320 -1575 4440 -1565
rect 4320 -1675 4330 -1575
rect 4430 -1675 4440 -1575
rect 4320 -1685 4440 -1675
rect 4320 -1905 4440 -1895
rect 4320 -2005 4330 -1905
rect 4430 -2005 4440 -1905
rect 4320 -2015 4440 -2005
rect 4320 -2235 4440 -2225
rect 4320 -2335 4330 -2235
rect 4430 -2335 4440 -2235
rect 4320 -2345 4440 -2335
rect 4320 -2565 4440 -2555
rect 4320 -2665 4330 -2565
rect 4430 -2665 4440 -2565
rect 4320 -2675 4440 -2665
rect 4320 -2895 4440 -2885
rect 4320 -2995 4330 -2895
rect 4430 -2995 4440 -2895
rect 4320 -3005 4440 -2995
rect 4320 -3225 4440 -3215
rect 4320 -3325 4330 -3225
rect 4430 -3325 4440 -3225
rect 4320 -3335 4440 -3325
rect 4320 -3555 4440 -3545
rect 4320 -3655 4330 -3555
rect 4430 -3655 4440 -3555
rect 4320 -3665 4440 -3655
rect 4320 -3885 4440 -3875
rect 4320 -3985 4330 -3885
rect 4430 -3985 4440 -3885
rect 4320 -3995 4440 -3985
rect 4320 -4215 4440 -4205
rect 4320 -4315 4330 -4215
rect 4430 -4315 4440 -4215
rect 4320 -4325 4440 -4315
rect 4320 -4545 4440 -4535
rect 4320 -4645 4330 -4545
rect 4430 -4645 4440 -4545
rect 4320 -4655 4440 -4645
rect 4320 -4875 4440 -4865
rect 4320 -4975 4330 -4875
rect 4430 -4975 4440 -4875
rect 4320 -4985 4440 -4975
rect 3900 -5205 4020 -5195
rect 3900 -5305 3910 -5205
rect 4010 -5305 4020 -5205
rect 3900 -5315 4020 -5305
rect 4320 -5205 4440 -5195
rect 4320 -5305 4330 -5205
rect 4430 -5305 4440 -5205
rect 4320 -5315 4440 -5305
<< via1 >>
rect 675 690 725 740
rect 2220 685 2270 735
rect 3730 680 3800 750
rect 4330 460 4430 560
rect 4330 -25 4430 75
rect 4330 -355 4430 -255
rect 4330 -685 4430 -585
rect 4330 -1015 4430 -915
rect 4330 -1345 4430 -1245
rect 4330 -1675 4430 -1575
rect 4330 -2005 4430 -1905
rect 4330 -2335 4430 -2235
rect 4330 -2665 4430 -2565
rect 4330 -2995 4430 -2895
rect 4330 -3325 4430 -3225
rect 4330 -3655 4430 -3555
rect 4330 -3985 4430 -3885
rect 4330 -4315 4430 -4215
rect 4330 -4645 4430 -4545
rect 4330 -4975 4430 -4875
rect 3910 -5305 4010 -5205
rect 4330 -5305 4430 -5205
<< metal2 >>
rect 3710 750 4120 775
rect 665 740 735 750
rect 665 690 675 740
rect 725 690 735 740
rect 665 680 735 690
rect 2210 735 2280 745
rect 2210 685 2220 735
rect 2270 685 2280 735
rect 2210 675 2280 685
rect 3710 680 3730 750
rect 3800 680 4120 750
rect 3710 655 4120 680
rect 4000 -3705 4120 655
rect 4325 560 4435 565
rect 4325 460 4330 560
rect 4430 460 4435 560
rect 4325 455 4435 460
rect 4320 75 4440 85
rect 4320 -25 4330 75
rect 4430 -25 4440 75
rect 4320 -35 4440 -25
rect 4320 -255 4440 -245
rect 4320 -355 4330 -255
rect 4430 -355 4440 -255
rect 4320 -365 4440 -355
rect 4320 -585 4440 -575
rect 4320 -685 4330 -585
rect 4430 -685 4440 -585
rect 4320 -695 4440 -685
rect 4320 -915 4440 -905
rect 4320 -1015 4330 -915
rect 4430 -1015 4440 -915
rect 4320 -1025 4440 -1015
rect 4320 -1245 4440 -1235
rect 4320 -1345 4330 -1245
rect 4430 -1345 4440 -1245
rect 4320 -1355 4440 -1345
rect 4320 -1575 4440 -1565
rect 4320 -1675 4330 -1575
rect 4430 -1675 4440 -1575
rect 4320 -1685 4440 -1675
rect 4320 -1905 4440 -1895
rect 4320 -2005 4330 -1905
rect 4430 -2005 4440 -1905
rect 4320 -2015 4440 -2005
rect 4320 -2235 4440 -2225
rect 4320 -2335 4330 -2235
rect 4430 -2335 4440 -2235
rect 4320 -2345 4440 -2335
rect 4320 -2565 4440 -2555
rect 4320 -2665 4330 -2565
rect 4430 -2665 4440 -2565
rect 4320 -2675 4440 -2665
rect 4320 -2895 4440 -2885
rect 4320 -2995 4330 -2895
rect 4430 -2995 4440 -2895
rect 4320 -3005 4440 -2995
rect 4320 -3225 4440 -3215
rect 4320 -3325 4330 -3225
rect 4430 -3325 4440 -3225
rect 4320 -3335 4440 -3325
rect 4320 -3555 4440 -3545
rect 4320 -3655 4330 -3555
rect 4430 -3655 4440 -3555
rect 4320 -3665 4440 -3655
rect 3458 -3715 4120 -3705
rect 3458 -3815 3468 -3715
rect 3568 -3815 4120 -3715
rect 3458 -3825 4120 -3815
rect 4320 -3885 4440 -3875
rect 4320 -3985 4330 -3885
rect 4430 -3985 4440 -3885
rect 4320 -3995 4440 -3985
rect 4320 -4215 4440 -4205
rect 4320 -4315 4330 -4215
rect 4430 -4315 4440 -4215
rect 4320 -4325 4440 -4315
rect 4320 -4545 4440 -4535
rect 4320 -4645 4330 -4545
rect 4430 -4645 4440 -4545
rect 4320 -4655 4440 -4645
rect 4320 -4875 4440 -4865
rect 4320 -4975 4330 -4875
rect 4430 -4975 4440 -4875
rect 4320 -4985 4440 -4975
rect 3900 -5205 4020 -5195
rect 3900 -5305 3910 -5205
rect 4010 -5305 4020 -5205
rect 3900 -5315 4020 -5305
rect 4320 -5205 4440 -5195
rect 4320 -5305 4330 -5205
rect 4430 -5305 4440 -5205
rect 4320 -5315 4440 -5305
<< via2 >>
rect 675 690 725 740
rect 2220 685 2270 735
rect 4330 460 4430 560
rect 4330 -25 4430 75
rect 4330 -355 4430 -255
rect 4330 -685 4430 -585
rect 4330 -1015 4430 -915
rect 4330 -1345 4430 -1245
rect 4330 -1675 4430 -1575
rect 4330 -2005 4430 -1905
rect 4330 -2335 4430 -2235
rect 4330 -2665 4430 -2565
rect 4330 -2995 4430 -2895
rect 4330 -3325 4430 -3225
rect 4330 -3655 4430 -3555
rect 3468 -3815 3568 -3715
rect 4330 -3985 4430 -3885
rect 4330 -4315 4430 -4215
rect 4330 -4645 4430 -4545
rect 4330 -4975 4430 -4875
rect 3910 -5305 4010 -5205
rect 4330 -5305 4430 -5205
<< metal3 >>
rect 665 740 735 750
rect 665 690 675 740
rect 725 690 735 740
rect 665 680 735 690
rect 2195 735 2295 760
rect 2195 685 2220 735
rect 2270 685 2295 735
rect 2195 210 2295 685
rect 4325 560 4435 565
rect 4325 460 4330 560
rect 4430 460 4435 560
rect 4325 455 4435 460
rect 2195 110 3890 210
rect 3790 -1920 3890 110
rect 4320 75 4440 85
rect 4320 -25 4330 75
rect 4430 -25 4440 75
rect 4320 -35 4440 -25
rect 4320 -255 4440 -245
rect 4320 -355 4330 -255
rect 4430 -355 4440 -255
rect 4320 -365 4440 -355
rect 4320 -585 4440 -575
rect 4320 -685 4330 -585
rect 4430 -685 4440 -585
rect 4320 -695 4440 -685
rect 4320 -915 4440 -905
rect 4320 -1015 4330 -915
rect 4430 -1015 4440 -915
rect 4320 -1025 4440 -1015
rect 4320 -1245 4440 -1235
rect 4320 -1345 4330 -1245
rect 4430 -1345 4440 -1245
rect 4320 -1355 4440 -1345
rect 4320 -1575 4440 -1565
rect 4320 -1675 4330 -1575
rect 4430 -1675 4440 -1575
rect 4320 -1685 4440 -1675
rect 3453 -1930 3890 -1920
rect 3453 -2030 3463 -1930
rect 3563 -2030 3890 -1930
rect 4320 -1905 4440 -1895
rect 4320 -2005 4330 -1905
rect 4430 -2005 4440 -1905
rect 4320 -2015 4440 -2005
rect 3453 -2040 3890 -2030
rect 4320 -2235 4440 -2225
rect 4320 -2335 4330 -2235
rect 4430 -2335 4440 -2235
rect 4320 -2345 4440 -2335
rect 4320 -2565 4440 -2555
rect 4320 -2665 4330 -2565
rect 4430 -2665 4440 -2565
rect 4320 -2675 4440 -2665
rect 4320 -2895 4440 -2885
rect 4320 -2995 4330 -2895
rect 4430 -2995 4440 -2895
rect 4320 -3005 4440 -2995
rect 4320 -3225 4440 -3215
rect 4320 -3325 4330 -3225
rect 4430 -3325 4440 -3225
rect 4320 -3335 4440 -3325
rect 4320 -3555 4440 -3545
rect 4320 -3655 4330 -3555
rect 4430 -3655 4440 -3555
rect 4320 -3665 4440 -3655
rect 3458 -3715 3578 -3705
rect 3458 -3815 3468 -3715
rect 3568 -3815 3578 -3715
rect 3458 -3825 3578 -3815
rect 4320 -3885 4440 -3875
rect 4320 -3985 4330 -3885
rect 4430 -3985 4440 -3885
rect 4320 -3995 4440 -3985
rect 4320 -4215 4440 -4205
rect 4320 -4315 4330 -4215
rect 4430 -4315 4440 -4215
rect 4320 -4325 4440 -4315
rect 4320 -4545 4440 -4535
rect 4320 -4645 4330 -4545
rect 4430 -4645 4440 -4545
rect 4320 -4655 4440 -4645
rect 4320 -4875 4440 -4865
rect 4320 -4975 4330 -4875
rect 4430 -4975 4440 -4875
rect 4320 -4985 4440 -4975
rect 3900 -5205 4020 -5195
rect 3900 -5305 3910 -5205
rect 4010 -5305 4020 -5205
rect 3900 -5315 4020 -5305
rect 4320 -5205 4440 -5195
rect 4320 -5305 4330 -5205
rect 4430 -5305 4440 -5205
rect 4320 -5315 4440 -5305
<< via3 >>
rect 675 690 725 740
rect 4330 460 4430 560
rect 4330 -25 4430 75
rect 4330 -355 4430 -255
rect 4330 -685 4430 -585
rect 4330 -1015 4430 -915
rect 4330 -1345 4430 -1245
rect 4330 -1675 4430 -1575
rect 3463 -2030 3563 -1930
rect 4330 -2005 4430 -1905
rect 4330 -2335 4430 -2235
rect 4330 -2665 4430 -2565
rect 4330 -2995 4430 -2895
rect 4330 -3325 4430 -3225
rect 4330 -3655 4430 -3555
rect 3468 -3815 3568 -3715
rect 4330 -3985 4430 -3885
rect 4330 -4315 4430 -4215
rect 4330 -4645 4430 -4545
rect 4330 -4975 4430 -4875
rect 3910 -5305 4010 -5205
rect 4330 -5305 4430 -5205
<< metal4 >>
rect 665 740 735 750
rect 665 690 675 740
rect 725 690 735 740
rect 665 680 735 690
rect 675 -205 725 680
rect 4305 560 4455 595
rect 4305 460 4330 560
rect 4430 460 4455 560
rect 4305 75 4455 460
rect 4305 -25 4330 75
rect 4430 -25 4455 75
rect 4305 -255 4455 -25
rect 4305 -355 4330 -255
rect 4430 -355 4455 -255
rect 4305 -585 4455 -355
rect 4305 -685 4330 -585
rect 4430 -685 4455 -585
rect 4305 -915 4455 -685
rect 4305 -1015 4330 -915
rect 4430 -1015 4455 -915
rect 4305 -1245 4455 -1015
rect 4305 -1345 4330 -1245
rect 4430 -1345 4455 -1245
rect 4305 -1575 4455 -1345
rect 4305 -1625 4330 -1575
rect 3965 -1675 4330 -1625
rect 4430 -1675 4455 -1575
rect 3965 -1775 4455 -1675
rect 4305 -1905 4455 -1775
rect 3453 -1930 3573 -1920
rect 3453 -2030 3463 -1930
rect 3563 -2030 3573 -1930
rect 3453 -2040 3573 -2030
rect 4305 -2005 4330 -1905
rect 4430 -2005 4455 -1905
rect 4305 -2235 4455 -2005
rect 4305 -2335 4330 -2235
rect 4430 -2335 4455 -2235
rect 4305 -2565 4455 -2335
rect 4305 -2665 4330 -2565
rect 4430 -2665 4455 -2565
rect 4305 -2895 4455 -2665
rect 4305 -2995 4330 -2895
rect 4430 -2995 4455 -2895
rect 4305 -3225 4455 -2995
rect 4305 -3325 4330 -3225
rect 4430 -3325 4455 -3225
rect 4305 -3395 4455 -3325
rect 3950 -3545 4455 -3395
rect 4305 -3555 4455 -3545
rect 4305 -3655 4330 -3555
rect 4430 -3655 4455 -3555
rect 3458 -3715 3578 -3705
rect 3458 -3815 3468 -3715
rect 3568 -3815 3578 -3715
rect 3458 -3825 3578 -3815
rect 4305 -3885 4455 -3655
rect 4305 -3985 4330 -3885
rect 4430 -3985 4455 -3885
rect 4305 -4215 4455 -3985
rect 4305 -4315 4330 -4215
rect 4430 -4315 4455 -4215
rect 4305 -4545 4455 -4315
rect 4305 -4645 4330 -4545
rect 4430 -4645 4455 -4545
rect 4305 -4875 4455 -4645
rect 4305 -4975 4330 -4875
rect 4430 -4975 4455 -4875
rect 4305 -5180 4455 -4975
rect 3885 -5205 4455 -5180
rect 3885 -5305 3910 -5205
rect 4010 -5305 4330 -5205
rect 4430 -5305 4455 -5205
rect 3885 -5330 4455 -5305
use cbank  cbank_1
timestamp 1647788355
transform 1 0 -42 0 1 -2705
box -15 -840 4075 775
use cbank  cbank_2
timestamp 1647788355
transform 1 0 -42 0 1 -4490
box -15 -840 4075 775
use cbank  cbank_0
timestamp 1647788355
transform 1 0 -42 0 1 -935
box -15 -840 4075 775
use ro_var_extend  ro_var_extend_0
timestamp 1640959680
transform 1 0 487 0 1 675
box -375 -595 3780 765
<< labels >>
rlabel locali 1123 -825 1123 -825 1 a0
rlabel locali 1617 -830 1617 -830 1 a1
rlabel locali 3673 -825 3673 -825 1 a5
rlabel locali 3072 -825 3072 -825 1 a4
rlabel locali 2591 -825 2591 -825 1 a3
rlabel locali 2101 -835 2101 -835 1 a2
rlabel space 3630 370 3630 370 1 vcont
rlabel space 1275 1115 1275 1115 1 vdd!
rlabel locali 3644 713 3644 713 1 out
<< end >>
