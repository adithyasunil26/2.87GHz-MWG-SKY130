magic
tech sky130A
timestamp 1711901915
<< checkpaint >>
rect 7639 2155 13908 10545
<< nwell >>
rect -3185 7805 -3090 9815
rect -3290 7585 -2985 7805
<< nsubdiff >>
rect -3210 7755 -3065 7770
rect -3210 7645 -3195 7755
rect -3080 7645 -3065 7755
rect -3210 7635 -3065 7645
<< nsubdiffcont >>
rect -3195 7645 -3080 7755
<< locali >>
rect -1502 10196 -1364 10217
rect -1502 10084 -1488 10196
rect -1378 10084 -1364 10196
rect -1502 10067 -1364 10084
rect -1499 9668 -1368 10067
rect 8310 9515 8778 9518
rect 7803 9114 8778 9515
rect 8310 9112 8778 9114
rect -5021 7604 -4961 7864
rect -3205 7755 -3070 7765
rect -3205 7645 -3195 7755
rect -3080 7645 -3070 7755
rect -3205 7640 -3070 7645
rect -5021 7545 -4477 7604
rect -4534 7380 -4479 7545
rect 7885 6690 8744 6954
rect -1492 6376 -1368 6388
rect -5053 5917 -4915 6349
rect -4015 5926 -3823 6332
rect -1492 6277 -1478 6376
rect -1382 6277 -1368 6376
rect -1492 6263 -1368 6277
rect -729 6145 82 6336
rect -2750 5215 -2700 5222
rect -2750 5179 -2743 5215
rect -2708 5179 -2700 5215
rect -2750 5139 -2700 5179
rect 7861 4862 8720 5126
rect -2265 4621 -2162 4628
rect -3003 4592 -2945 4595
rect -2265 4592 -2254 4621
rect -3003 4590 -2788 4592
rect -3003 4547 -2994 4590
rect -2951 4552 -2788 4590
rect -2951 4550 -2906 4552
rect -2606 4550 -2254 4592
rect -2951 4547 -2945 4550
rect -2320 4549 -2254 4550
rect -3003 4538 -2945 4547
rect -2265 4529 -2254 4549
rect -2170 4529 -2162 4621
rect -2265 4525 -2162 4529
rect -4902 4072 -4702 4384
rect -4254 4037 -3882 4394
rect -3547 4326 -2730 4356
rect -331 3685 129 3956
rect -378 2878 294 3207
rect 7919 3059 8768 3323
rect -331 2025 129 2296
<< viali >>
rect -1488 10084 -1378 10196
rect 9501 9577 9574 9642
rect -3195 7645 -3080 7755
rect -1478 6277 -1382 6376
rect -2743 5179 -2708 5215
rect -2994 4547 -2951 4590
rect -2254 4529 -2170 4621
rect -515 2395 -490 2420
<< metal1 >>
rect -1502 10196 -1364 10217
rect -1502 10084 -1488 10196
rect -1378 10084 -1364 10196
rect -1502 10067 -1364 10084
rect 9485 9642 9591 9654
rect 9485 9577 9501 9642
rect 9574 9577 9591 9642
rect 9485 9566 9591 9577
rect 3986 9380 4062 9382
rect 380 9370 4062 9380
rect 380 9245 8140 9370
rect -3205 7755 -3070 7765
rect -3205 7645 -3195 7755
rect -3080 7645 -3070 7755
rect -3205 7640 -3070 7645
rect 380 7630 460 9245
rect 8065 8900 8140 9245
rect 8065 8899 8575 8900
rect 8065 8810 9181 8899
rect 8065 8805 8140 8810
rect 8526 8805 9181 8810
rect -595 7510 465 7630
rect 380 7505 460 7510
rect -1492 6376 -1368 6388
rect -1492 6277 -1478 6376
rect -1382 6277 -1368 6376
rect -1492 6263 -1368 6277
rect -3354 5530 -3086 5534
rect -3375 5515 -3086 5530
rect -3354 5503 -3086 5515
rect -3320 5405 -3275 5410
rect -3320 5395 -3315 5405
rect -3375 5380 -3315 5395
rect -3320 5370 -3315 5380
rect -3280 5370 -3275 5405
rect -3320 5365 -3275 5370
rect -3119 4576 -3086 5503
rect -2750 5215 -2700 5222
rect -2750 5179 -2743 5215
rect -2708 5179 -2700 5215
rect -2750 5170 -2700 5179
rect -2265 4621 -2162 4628
rect -3003 4590 -2945 4595
rect -3003 4576 -2994 4590
rect -3122 4550 -2994 4576
rect -3003 4547 -2994 4550
rect -2951 4547 -2945 4590
rect -3003 4538 -2945 4547
rect -2265 4529 -2254 4621
rect -2170 4529 -2162 4621
rect -2265 4525 -2162 4529
rect -525 2425 -480 2430
rect -525 2390 -520 2425
rect -485 2390 -480 2425
rect -525 2385 -480 2390
<< via1 >>
rect -1488 10084 -1378 10196
rect 9501 9577 9574 9642
rect -3195 7645 -3080 7755
rect -1478 6277 -1382 6376
rect -3315 5370 -3280 5405
rect -2743 5179 -2708 5215
rect -2254 4529 -2170 4621
rect -520 2420 -485 2425
rect -520 2395 -515 2420
rect -515 2395 -490 2420
rect -490 2395 -485 2420
rect -520 2390 -485 2395
<< metal2 >>
rect -74 10223 -50 10224
rect -74 10222 129 10223
rect -1502 10196 129 10222
rect -1502 10084 -1488 10196
rect -1378 10084 129 10196
rect -1502 10067 129 10084
rect -110 10063 129 10067
rect -61 8322 129 10063
rect 9485 9642 9591 9654
rect 9485 9577 9501 9642
rect 9574 9577 9591 9642
rect 9485 9566 9591 9577
rect -3205 7755 -3070 7765
rect -3205 7645 -3195 7755
rect -3080 7645 -3070 7755
rect -3205 7640 -3070 7645
rect -67 7397 129 8322
rect -73 7340 129 7397
rect -1492 6376 -1368 6388
rect -1492 6277 -1478 6376
rect -1382 6277 -1368 6376
rect -1492 6263 -1368 6277
rect -73 6071 127 7340
rect -5100 5575 -4960 5590
rect -3325 5405 -3270 5415
rect -3325 5370 -3315 5405
rect -3280 5370 -3270 5405
rect -3325 5360 -3270 5370
rect -2750 5215 -2700 5222
rect -2750 5179 -2743 5215
rect -2708 5179 -2700 5215
rect -2750 5170 -2700 5179
rect -5250 4720 -4960 4740
rect -5250 1991 -5200 4720
rect -79 4623 130 6071
rect -2264 4621 130 4623
rect -2264 4529 -2254 4621
rect -2170 4529 130 4621
rect -2264 4523 130 4529
rect -79 4518 130 4523
rect 12610 4220 12740 4935
rect -5160 4185 12740 4220
rect -5160 2435 -5140 4185
rect -4675 3800 -4625 3810
rect -4675 3770 -4665 3800
rect -4635 3770 -4625 3800
rect -4675 3760 -4625 3770
rect -5160 2415 -5095 2435
rect -530 2425 -475 2435
rect -530 2390 -520 2425
rect -485 2390 -475 2425
rect -530 2380 -475 2390
rect -5250 1990 -5096 1991
rect -525 1990 -490 2380
rect -5250 1950 -490 1990
rect -5250 1949 -5200 1950
rect -5165 1949 -5135 1950
<< via2 >>
rect 9501 9577 9574 9642
rect -3195 7645 -3080 7755
rect -1478 6277 -1382 6376
rect -3315 5370 -3280 5405
rect -2743 5179 -2708 5215
rect -4665 3770 -4635 3800
<< metal3 >>
rect 9485 9642 9591 9654
rect 9485 9577 9501 9642
rect 9574 9577 9591 9642
rect 9485 9566 9591 9577
rect -3290 7755 -2985 7805
rect -3290 7645 -3195 7755
rect -3080 7645 -2985 7755
rect -3290 7585 -2985 7645
rect -1500 6376 -1349 6388
rect -1500 6277 -1478 6376
rect -1382 6277 -1349 6376
rect -3331 5431 -2069 5433
rect -1500 5431 -1349 6277
rect -3331 5405 -1349 5431
rect -3331 5370 -3315 5405
rect -3280 5370 -1349 5405
rect -3331 5346 -1349 5370
rect -1500 5339 -1349 5346
rect -2750 5215 -2700 5222
rect -2750 5179 -2743 5215
rect -2708 5179 -2700 5215
rect -2750 5170 -2700 5179
rect -4675 3805 -4625 3810
rect -4675 3765 -4670 3805
rect -4630 3765 -4625 3805
rect -4675 3760 -4625 3765
<< via3 >>
rect 9501 9577 9574 9642
rect -3195 7645 -3080 7755
rect -2743 5179 -2708 5215
rect -4670 3800 -4630 3805
rect -4670 3770 -4665 3800
rect -4665 3770 -4635 3800
rect -4635 3770 -4630 3800
rect -4670 3765 -4630 3770
<< metal4 >>
rect 9339 10823 9609 10829
rect -92 10814 9609 10823
rect -3926 10808 9609 10814
rect -5794 10779 -5174 10780
rect -4316 10779 9609 10808
rect -5794 10552 9609 10779
rect -5794 10510 -3711 10552
rect -92 10543 9609 10552
rect 9339 10541 9609 10543
rect -5794 10509 -4166 10510
rect -5794 10504 -5174 10509
rect -5790 5810 -5439 10504
rect -3896 10488 -3715 10510
rect -3895 10110 -3716 10488
rect -3898 10099 -3716 10110
rect -3898 9708 -3719 10099
rect -3185 7780 -3090 9815
rect 9470 9642 9607 10541
rect 9470 9577 9501 9642
rect 9574 9577 9607 9642
rect 9470 9552 9607 9577
rect -3210 7755 -3055 7780
rect -3210 7645 -3195 7755
rect -3080 7645 -3055 7755
rect -3210 7625 -3055 7645
rect -5790 5720 -4891 5810
rect -2751 5757 -2701 5758
rect -3387 5727 -2701 5757
rect -5790 3871 -5439 5720
rect -3377 5654 -3293 5727
rect -2751 5222 -2701 5727
rect -2751 5215 -2700 5222
rect -2751 5179 -2743 5215
rect -2708 5179 -2700 5215
rect -2751 5170 -2700 5179
rect -2751 5164 -2701 5170
rect -4660 3897 -4595 3900
rect -4769 3871 -4595 3897
rect -5790 3860 -4595 3871
rect -5790 3845 -4625 3860
rect -5790 3826 -4716 3845
rect -5790 3260 -5439 3826
rect -4659 3814 -4625 3845
rect -4660 3810 -4625 3814
rect -4675 3805 -4625 3810
rect -4675 3765 -4670 3805
rect -4630 3765 -4625 3805
rect -4675 3760 -4625 3765
rect -5791 3090 -4643 3260
use ro_complete  ro_complete_0
timestamp 1647788355
transform 1 0 8617 0 1 8475
box -348 -5690 4661 1440
use inverter  inverter_0
timestamp 1647877520
transform 1 0 -2894 0 1 4593
box 75 -311 310 557
use cp  cp_0
timestamp 1640911461
transform 1 0 -4895 0 1 7840
box -415 -1715 4690 2035
use filter  filter_0
timestamp 1640983258
transform 1 0 1810 0 1 10450
box -1800 -11005 6240 390
use divider  divider_0
timestamp 1647769399
transform 1 0 -4910 0 1 1985
box -490 -235 4690 2150
use pd  pd_0
timestamp 1711730514
transform 1 0 -4845 0 1 5180
box -215 -855 1685 810
<< labels >>
rlabel locali -3140 7755 -3140 7755 1 vdd!
rlabel metal4 -3755 9794 -3755 9795 1 vdd!
rlabel metal2 -4810 1956 -4810 1956 1 div
rlabel metal2 -2696 4201 -2696 4201 1 vco
rlabel metal2 -5084 5583 -5084 5583 1 ref
rlabel locali -74 3770 -74 3770 1 gnd!
rlabel space 9739 6638 9739 6638 1 a0
rlabel space 10231 6623 10231 6623 1 a1
rlabel space 10721 6626 10721 6626 1 a2
rlabel space 11204 6625 11204 6625 1 a3
rlabel space 11694 6604 11694 6604 1 a4
rlabel space 12292 6623 12292 6623 1 a5
<< end >>
