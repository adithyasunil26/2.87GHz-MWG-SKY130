magic
tech sky130A
magscale 1 2
timestamp 1712611811
<< ndiff >>
rect 1720 -30 1860 110
rect 2730 92 2870 110
rect 2730 -8 2750 92
rect 2850 -8 2870 92
rect 2730 -30 2870 -8
rect 3680 92 3820 110
rect 3680 -8 3700 92
rect 3800 -8 3820 92
rect 3680 -30 3820 -8
rect 4660 92 4800 110
rect 4660 -8 4680 92
rect 4780 -8 4800 92
rect 4660 -30 4800 -8
rect 5640 92 5780 110
rect 5640 -8 5660 92
rect 5760 -8 5780 92
rect 5640 -30 5780 -8
rect 6660 92 6800 110
rect 6660 -8 6680 92
rect 6780 -8 6800 92
rect 6660 -30 6800 -8
<< ndiffc >>
rect 2750 -8 2850 92
rect 3700 -8 3800 92
rect 4680 -8 4780 92
rect 5660 -8 5760 92
rect 6680 -8 6780 92
<< psubdiff >>
rect 950 -1430 1210 -1400
rect 950 -1630 980 -1430
rect 1180 -1630 1210 -1430
rect 950 -1660 1210 -1630
rect 4850 -1430 5110 -1400
rect 4850 -1630 4880 -1430
rect 5080 -1630 5110 -1430
rect 4850 -1660 5110 -1630
<< psubdiffcont >>
rect 980 -1630 1180 -1430
rect 4880 -1630 5080 -1430
<< locali >>
rect 1000 1360 1190 1380
rect 1000 1230 1020 1360
rect 970 1210 1020 1230
rect 1170 1210 1190 1360
rect 970 1190 1190 1210
rect 1990 190 2000 260
rect 3000 190 3010 260
rect 3950 190 3960 260
rect 4930 190 4940 260
rect 5910 190 5920 260
rect 6930 190 6940 260
rect 1720 90 1860 110
rect 1720 -10 1740 90
rect 1840 -10 1860 90
rect 1720 -30 1860 -10
rect 2730 92 2870 110
rect 2730 -10 2750 92
rect 2850 -10 2870 92
rect 2730 -30 2870 -10
rect 3680 92 3820 110
rect 3680 -10 3700 92
rect 3800 -10 3820 92
rect 3680 -30 3820 -10
rect 4660 92 4800 110
rect 4660 -10 4680 92
rect 4780 -10 4800 92
rect 4660 -30 4800 -10
rect 5640 92 5780 110
rect 5640 -10 5660 92
rect 5760 -10 5780 92
rect 5640 -30 5780 -10
rect 6660 92 6800 110
rect 6660 -10 6680 92
rect 6780 -10 6800 92
rect 6660 -30 6800 -10
rect 1990 -1410 2090 -1270
rect 3000 -1410 3100 -1280
rect 3950 -1410 4050 -1280
rect 4930 -1410 5030 -1280
rect 5910 -1410 6010 -1280
rect 6930 -1410 7030 -1280
rect 960 -1430 1200 -1410
rect 960 -1630 980 -1430
rect 1180 -1630 1200 -1430
rect 960 -1650 1200 -1630
rect 1920 -1430 2160 -1410
rect 1920 -1630 1940 -1430
rect 2140 -1630 2160 -1430
rect 1920 -1650 2160 -1630
rect 2930 -1430 3170 -1410
rect 2930 -1630 2950 -1430
rect 3150 -1630 3170 -1430
rect 2930 -1650 3170 -1630
rect 3880 -1430 4120 -1410
rect 3880 -1630 3900 -1430
rect 4100 -1630 4120 -1430
rect 3880 -1650 4120 -1630
rect 4860 -1430 5100 -1410
rect 4860 -1630 4880 -1430
rect 5080 -1630 5100 -1430
rect 4860 -1650 5100 -1630
rect 5840 -1430 6080 -1410
rect 5840 -1630 5860 -1430
rect 6060 -1630 6080 -1430
rect 5840 -1650 6080 -1630
rect 6870 -1430 7110 -1410
rect 6870 -1630 6890 -1430
rect 7090 -1630 7110 -1430
rect 6870 -1650 7110 -1630
<< viali >>
rect 1020 1210 1170 1360
rect 1740 -10 1840 90
rect 2750 -8 2850 90
rect 2750 -10 2850 -8
rect 3700 -8 3800 90
rect 3700 -10 3800 -8
rect 4680 -8 4780 90
rect 4680 -10 4780 -8
rect 5660 -8 5760 90
rect 5660 -10 5760 -8
rect 6680 -8 6780 90
rect 6680 -10 6780 -8
rect 980 -1630 1180 -1430
rect 1940 -1630 2140 -1430
rect 2950 -1630 3150 -1430
rect 3900 -1630 4100 -1430
rect 4880 -1630 5080 -1430
rect 5860 -1630 6060 -1430
rect 6890 -1630 7090 -1430
<< metal1 >>
rect 1000 1360 1190 1380
rect 1000 1210 1020 1360
rect 1170 1210 1190 1360
rect 1000 1190 1190 1210
rect 1720 90 1860 110
rect 1720 -10 1740 90
rect 1840 -10 1860 90
rect 1720 -30 1860 -10
rect 2730 90 2870 110
rect 2730 -10 2750 90
rect 2850 -10 2870 90
rect 2730 -30 2870 -10
rect 3680 90 3820 110
rect 3680 -10 3700 90
rect 3800 -10 3820 90
rect 3680 -30 3820 -10
rect 4660 90 4800 110
rect 4660 -10 4680 90
rect 4780 -10 4800 90
rect 4660 -30 4800 -10
rect 5640 90 5780 110
rect 5640 -10 5660 90
rect 5760 -10 5780 90
rect 5640 -30 5780 -10
rect 6660 90 6800 110
rect 6660 -10 6680 90
rect 6780 -10 6800 90
rect 6660 -30 6800 -10
rect 960 -1430 1200 -1410
rect 960 -1630 980 -1430
rect 1180 -1630 1200 -1430
rect 960 -1650 1200 -1630
rect 1920 -1430 2160 -1410
rect 1920 -1630 1940 -1430
rect 2140 -1630 2160 -1430
rect 1920 -1650 2160 -1630
rect 2930 -1430 3170 -1410
rect 2930 -1630 2950 -1430
rect 3150 -1630 3170 -1430
rect 2930 -1650 3170 -1630
rect 3880 -1430 4120 -1410
rect 3880 -1630 3900 -1430
rect 4100 -1630 4120 -1430
rect 3880 -1650 4120 -1630
rect 4860 -1430 5100 -1410
rect 4860 -1630 4880 -1430
rect 5080 -1630 5100 -1430
rect 4860 -1650 5100 -1630
rect 5840 -1430 6080 -1410
rect 5840 -1630 5860 -1430
rect 6060 -1630 6080 -1430
rect 5840 -1650 6080 -1630
rect 6870 -1430 7110 -1410
rect 6870 -1630 6890 -1430
rect 7090 -1630 7110 -1430
rect 6870 -1650 7110 -1630
<< via1 >>
rect 1020 1210 1170 1360
rect 1740 -10 1840 90
rect 2750 -10 2850 90
rect 3700 -10 3800 90
rect 4680 -10 4780 90
rect 5660 -10 5760 90
rect 6680 -10 6780 90
rect 980 -1630 1180 -1430
rect 1940 -1630 2140 -1430
rect 2950 -1630 3150 -1430
rect 3900 -1630 4100 -1430
rect 4880 -1630 5080 -1430
rect 5860 -1630 6060 -1430
rect 6890 -1630 7090 -1430
<< metal2 >>
rect 1000 1360 1190 1380
rect 1000 1210 1020 1360
rect 1170 1210 1190 1360
rect 1000 1190 1190 1210
rect 1720 90 1860 110
rect 1720 -10 1740 90
rect 1840 -10 1860 90
rect 1720 -30 1860 -10
rect 2730 90 2870 110
rect 2730 -10 2750 90
rect 2850 -10 2870 90
rect 2730 -30 2870 -10
rect 3680 90 3820 110
rect 3680 -10 3700 90
rect 3800 -10 3820 90
rect 3680 -30 3820 -10
rect 4660 90 4800 110
rect 4660 -10 4680 90
rect 4780 -10 4800 90
rect 4660 -30 4800 -10
rect 5640 90 5780 110
rect 5640 -10 5660 90
rect 5760 -10 5780 90
rect 5640 -30 5780 -10
rect 6660 90 6800 110
rect 6660 -10 6680 90
rect 6780 -10 6800 90
rect 6660 -30 6800 -10
rect 960 -1430 1200 -1410
rect 960 -1630 980 -1430
rect 1180 -1630 1200 -1430
rect 960 -1650 1200 -1630
rect 1920 -1430 2160 -1410
rect 1920 -1630 1940 -1430
rect 2140 -1630 2160 -1430
rect 1920 -1650 2160 -1630
rect 2930 -1430 3170 -1410
rect 2930 -1630 2950 -1430
rect 3150 -1630 3170 -1430
rect 2930 -1650 3170 -1630
rect 3880 -1430 4120 -1410
rect 3880 -1630 3900 -1430
rect 4100 -1630 4120 -1430
rect 3880 -1650 4120 -1630
rect 4860 -1430 5100 -1410
rect 4860 -1630 4880 -1430
rect 5080 -1630 5100 -1430
rect 4860 -1650 5100 -1630
rect 5840 -1430 6080 -1410
rect 5840 -1630 5860 -1430
rect 6060 -1630 6080 -1430
rect 5840 -1650 6080 -1630
rect 6870 -1430 7110 -1410
rect 6870 -1630 6890 -1430
rect 7090 -1630 7110 -1430
rect 6870 -1650 7110 -1630
<< via2 >>
rect 1020 1210 1170 1360
rect 1740 -10 1840 90
rect 2750 -10 2850 90
rect 3700 -10 3800 90
rect 4680 -10 4780 90
rect 5660 -10 5760 90
rect 6680 -10 6780 90
rect 980 -1630 1180 -1430
rect 1940 -1630 2140 -1430
rect 2950 -1630 3150 -1430
rect 3900 -1630 4100 -1430
rect 4880 -1630 5080 -1430
rect 5860 -1630 6060 -1430
rect 6890 -1630 7090 -1430
<< metal3 >>
rect 1000 1360 1190 1380
rect 1000 1210 1020 1360
rect 1170 1210 1190 1360
rect 1000 1190 1190 1210
rect 1450 490 2200 1090
rect 2440 490 3190 1090
rect 3430 490 4180 1090
rect 4420 490 5170 1090
rect 5410 490 6160 1090
rect 6410 490 7160 1090
rect 1720 90 1860 490
rect 1720 -10 1740 90
rect 1840 -10 1860 90
rect 1720 -30 1860 -10
rect 2730 90 2870 490
rect 2730 -10 2750 90
rect 2850 -10 2870 90
rect 2730 -30 2870 -10
rect 3680 90 3820 490
rect 3680 -10 3700 90
rect 3800 -10 3820 90
rect 3680 -30 3820 -10
rect 4660 90 4800 490
rect 4660 -10 4680 90
rect 4780 -10 4800 90
rect 4660 -30 4800 -10
rect 5640 90 5780 490
rect 5640 -10 5660 90
rect 5760 -10 5780 90
rect 5640 -30 5780 -10
rect 6660 90 6800 490
rect 6660 -10 6680 90
rect 6780 -10 6800 90
rect 6660 -30 6800 -10
rect 960 -1430 1200 -1410
rect 960 -1630 980 -1430
rect 1180 -1630 1200 -1430
rect 960 -1650 1200 -1630
rect 1920 -1430 2160 -1410
rect 1920 -1630 1940 -1430
rect 2140 -1630 2160 -1430
rect 1920 -1650 2160 -1630
rect 2930 -1430 3170 -1410
rect 2930 -1630 2950 -1430
rect 3150 -1630 3170 -1430
rect 2930 -1650 3170 -1630
rect 3880 -1430 4120 -1410
rect 3880 -1630 3900 -1430
rect 4100 -1630 4120 -1430
rect 3880 -1650 4120 -1630
rect 4860 -1430 5100 -1410
rect 4860 -1630 4880 -1430
rect 5080 -1630 5100 -1430
rect 4860 -1650 5100 -1630
rect 5840 -1430 6080 -1410
rect 5840 -1630 5860 -1430
rect 6060 -1630 6080 -1430
rect 5840 -1650 6080 -1630
rect 6870 -1430 7110 -1410
rect 6870 -1630 6890 -1430
rect 7090 -1630 7110 -1430
rect 6870 -1650 7110 -1630
<< via3 >>
rect 1020 1210 1170 1360
rect 980 -1630 1180 -1430
rect 1940 -1630 2140 -1430
rect 2950 -1630 3150 -1430
rect 3900 -1630 4100 -1430
rect 4880 -1630 5080 -1430
rect 5860 -1630 6060 -1430
rect 6890 -1630 7090 -1430
<< mimcap >>
rect 1550 950 2110 990
rect 1550 630 1590 950
rect 2070 630 2110 950
rect 1550 590 2110 630
rect 2540 950 3100 990
rect 2540 630 2580 950
rect 3060 630 3100 950
rect 2540 590 3100 630
rect 3530 950 4090 990
rect 3530 630 3570 950
rect 4050 630 4090 950
rect 3530 590 4090 630
rect 4520 950 5080 990
rect 4520 630 4560 950
rect 5040 630 5080 950
rect 4520 590 5080 630
rect 5510 950 6070 990
rect 5510 630 5550 950
rect 6030 630 6070 950
rect 5510 590 6070 630
rect 6510 950 7070 990
rect 6510 630 6550 950
rect 7030 630 7070 950
rect 6510 590 7070 630
<< mimcapcontact >>
rect 1590 630 2070 950
rect 2580 630 3060 950
rect 3570 630 4050 950
rect 4560 630 5040 950
rect 5550 630 6030 950
rect 6550 630 7030 950
<< metal4 >>
rect 990 1360 7220 1390
rect 990 1210 1020 1360
rect 1170 1210 7220 1360
rect 990 1180 7220 1210
rect 1690 951 1890 1180
rect 2680 951 2880 1180
rect 3670 951 3870 1180
rect 4660 951 4860 1180
rect 5650 951 5850 1180
rect 6650 951 6850 1180
rect 1589 950 2071 951
rect 1589 630 1590 950
rect 2070 630 2071 950
rect 1589 629 2071 630
rect 2579 950 3061 951
rect 2579 630 2580 950
rect 3060 630 3061 950
rect 2579 629 3061 630
rect 3569 950 4051 951
rect 3569 630 3570 950
rect 4050 630 4051 950
rect 3569 629 4051 630
rect 4559 950 5041 951
rect 4559 630 4560 950
rect 5040 630 5041 950
rect 4559 629 5041 630
rect 5549 950 6031 951
rect 5549 630 5550 950
rect 6030 630 6031 950
rect 5549 629 6031 630
rect 6549 950 7031 951
rect 6549 630 6550 950
rect 7030 630 7031 950
rect 6549 629 7031 630
rect 930 -1380 1230 -242
rect 930 -1430 8150 -1380
rect 930 -1630 980 -1430
rect 1180 -1630 1940 -1430
rect 2140 -1630 2950 -1430
rect 3150 -1630 3900 -1430
rect 4100 -1630 4880 -1430
rect 5080 -1630 5860 -1430
rect 6060 -1630 6890 -1430
rect 7090 -1630 8150 -1430
rect 930 -1680 8150 -1630
use switch  switch_5
timestamp 1640608635
transform 1 0 6830 0 1 -1308
box -190 -40 240 1600
use switch  switch_4
timestamp 1640608635
transform 1 0 5810 0 1 -1308
box -190 -40 240 1600
use switch  switch_3
timestamp 1640608635
transform 1 0 4830 0 1 -1308
box -190 -40 240 1600
use switch  switch_2
timestamp 1640608635
transform 1 0 3850 0 1 -1308
box -190 -40 240 1600
use switch  switch_1
timestamp 1640608635
transform 1 0 2900 0 1 -1308
box -190 -40 240 1600
use switch  switch_0
timestamp 1640608635
transform 1 0 1890 0 1 -1308
box -190 -40 240 1600
<< labels >>
rlabel locali 2000 220 2000 220 1 a0
rlabel locali 3010 220 3010 220 1 a1
rlabel locali 3960 210 3960 210 1 a2
rlabel locali 4950 -1370 4951 -1370 1 gnd!
rlabel locali 4940 210 4940 210 1 a3
rlabel locali 5920 200 5920 200 1 a4
rlabel locali 6940 200 6940 200 1 a5
rlabel locali 980 1200 980 1200 1 v
<< end >>
