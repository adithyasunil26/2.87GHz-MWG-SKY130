* SPICE3 file created from ro_complete_buffered.ext - technology: sky130A

.lib "<path_to_pdk>/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

.global vdd gnd
Vdd vdd gnd 1.8

* Va0 a0 gnd pwl(0 0 9n 0 10n 1.8 100n 1.8)
* Va1 a1 gnd pwl(0 0 19n 0 20n 1.8 100n 1.8)
* Va2 a2 gnd pwl(0 0 29n 0 30n 1.8 100n 1.8)
* Va3 a3 gnd pwl(0 0 39n 0 40n 1.8 100n 1.8)
* Va4 a4 gnd pwl(0 0 49n 0 50n 1.8 100n 1.8)
* Va5 a5 gnd pwl(0 0 59n 0 60n 1.8 100n 1.8)
Va0 a0 gnd 0
Va1 a1 gnd 0
Va2 a2 gnd 0
Va3 a3 gnd 0
Va4 a4 gnd 0
Va5 a5 gnd 0
Vcont vcont gnd pwl(0 0 100n 1.8)

X0 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X14 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X17 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X26 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X30 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X34 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X35 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X40 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X43 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X49 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X60 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X61 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X64 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X65 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X72 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X76 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X80 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X82 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X85 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X87 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X88 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X90 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X91 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X93 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X94 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X95 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X97 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X98 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X100 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X102 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X103 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X104 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X105 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X106 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X107 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X108 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X109 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X110 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X111 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X112 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X113 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X115 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X117 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X119 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X120 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X121 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X122 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X123 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X124 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X125 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X126 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X127 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X128 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X129 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X130 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X131 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X132 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X133 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X134 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X136 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X137 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X138 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X139 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X141 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X142 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X143 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X144 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X145 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X146 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X147 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X148 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X149 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X150 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X151 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X152 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X153 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X154 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X157 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X158 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X159 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X160 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X161 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X162 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X163 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X164 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X165 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X166 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X167 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X168 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X169 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X170 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X171 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X172 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X173 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X174 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X175 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X176 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X177 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X178 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X179 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X180 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X181 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X182 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X183 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X184 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X185 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X186 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X187 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X188 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X189 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X190 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X191 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X192 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X193 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X194 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X195 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X196 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X197 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X198 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X199 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X200 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X201 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X202 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X203 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X204 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X205 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X206 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X207 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X208 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X209 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X210 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X211 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X212 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X213 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X214 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X215 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X216 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X217 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X218 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X219 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X220 tapered_buf_2/a_160_230# tapered_buf_2/in tapered_buf_2/a_n10_230# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X221 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X222 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X223 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X224 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X225 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X226 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X227 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X228 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X229 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X230 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X231 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X232 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X234 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X235 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X236 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X237 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X238 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X239 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X240 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X241 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X243 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X244 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X245 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X246 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X247 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X248 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X249 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X250 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X251 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X252 tapered_buf_2/a_580_0# tapered_buf_2/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X253 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X254 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X255 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X256 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X257 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X258 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X259 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X260 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X261 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X262 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X263 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X264 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X265 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X266 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X267 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X268 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X269 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X271 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X272 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X273 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X274 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X275 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X276 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X277 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X279 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X280 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X281 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X282 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X283 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X284 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X285 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X286 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X287 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X288 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X289 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X290 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X291 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X292 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X293 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X294 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X295 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X296 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X297 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X298 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X299 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X300 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X301 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X302 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X303 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X304 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X305 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X306 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X307 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X308 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X309 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X310 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X311 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X312 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X313 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X314 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X315 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X316 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X317 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X318 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X319 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X320 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X321 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X322 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X323 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X324 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X325 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X326 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X327 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X328 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X329 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X330 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X331 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X332 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X333 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X334 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X335 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X336 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X337 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X338 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X339 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X340 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X341 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X342 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X343 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X344 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X345 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X346 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X347 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X348 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X349 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X350 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X351 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X352 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X353 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X354 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X355 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X356 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X357 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X358 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X359 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X360 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X361 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X362 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X363 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X364 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X365 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X366 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X367 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X368 gnd tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X369 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X370 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X371 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X372 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X373 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X374 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X375 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X376 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X377 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X378 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X379 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X380 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X381 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X382 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X383 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X384 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X385 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X386 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X387 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X388 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X389 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X390 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X391 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X392 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X393 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X394 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X395 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X396 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X397 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X398 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X399 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X400 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X401 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X402 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X403 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X404 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X405 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X406 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X407 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X408 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X409 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X410 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X411 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X412 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X413 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X414 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X415 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X416 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X417 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X418 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X419 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X420 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X421 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X422 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X423 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X424 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X425 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X426 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X427 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X428 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X429 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X430 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X431 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X432 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X433 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X434 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X435 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X436 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X437 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X438 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X439 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X440 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X441 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X442 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X443 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X444 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X445 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X446 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X447 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X448 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X449 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X450 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X451 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X452 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X453 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X454 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X455 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X456 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X457 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X458 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X459 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X460 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X461 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X462 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X463 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X464 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X465 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X466 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X467 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X468 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X469 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X470 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X471 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X472 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X473 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X474 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X475 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X476 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X477 gnd tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X478 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X479 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X480 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X481 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X482 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X483 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X484 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X485 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X486 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X487 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X488 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X489 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X490 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X491 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X492 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X493 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X494 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X495 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X496 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X497 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X498 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X499 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X500 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X501 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X502 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X503 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X504 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X505 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X506 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X507 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X508 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X509 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X510 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X511 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X512 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X513 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X514 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X515 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X516 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X517 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X518 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X519 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X520 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X521 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X522 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X523 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X524 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X525 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X526 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X527 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X528 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X529 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X530 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X531 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X532 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X533 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X534 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X535 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X536 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X537 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X538 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X539 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X540 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X541 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X542 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X543 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X544 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X545 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X546 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X547 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X548 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X549 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X550 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X551 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X552 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X553 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X554 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X555 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X556 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X557 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X558 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X559 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X560 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X561 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X562 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X563 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X564 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X565 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X566 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X567 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X568 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X569 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X570 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X571 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X572 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X573 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X574 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X575 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X576 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X577 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X578 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X579 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X580 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X581 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X582 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X583 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X584 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X585 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X586 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X587 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X588 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X589 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X590 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X591 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X592 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X593 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X594 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X595 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X596 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X597 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X598 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X599 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X600 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X601 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X602 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X603 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X604 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X605 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X606 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X607 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X608 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X609 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X610 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X611 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X612 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X613 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X614 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X615 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X616 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X617 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X618 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X619 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X620 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X621 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X622 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X623 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X624 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X625 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X626 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X627 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X628 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X629 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X630 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X631 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X632 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X633 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X634 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X635 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X636 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X637 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X638 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X639 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X640 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X641 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X642 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X643 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X644 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X645 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X646 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X647 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X648 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X649 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X650 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X651 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X652 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X653 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X654 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X655 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X656 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X657 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X658 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X659 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X660 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X661 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X662 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X663 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X664 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X665 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X666 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X667 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X668 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X669 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X670 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X671 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X672 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X673 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X674 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X675 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X676 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X677 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X678 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X679 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X680 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X681 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X682 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X683 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X684 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X685 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X686 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X687 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X688 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X689 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X690 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X691 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X692 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X693 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X694 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X695 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X696 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X697 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X698 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X699 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X700 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X701 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X702 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X703 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X704 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X705 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X706 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X707 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X708 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X709 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X710 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X711 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X712 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X713 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X714 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X715 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X716 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X717 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X718 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X719 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X720 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X721 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X722 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X723 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X724 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X725 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X726 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X727 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X728 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X729 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X730 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X731 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X732 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X733 tapered_buf_2/a_580_0# tapered_buf_2/a_160_n140# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X734 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X735 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X736 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X737 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X738 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X739 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X740 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X741 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X742 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X743 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X744 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X745 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X746 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X747 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X748 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X749 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X750 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X751 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X752 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X753 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X754 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X755 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X756 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X757 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X758 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X759 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X760 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X761 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X762 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X763 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X764 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X765 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X766 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X767 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X768 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X769 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X770 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X771 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X772 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X773 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X774 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X775 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X776 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X777 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X778 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X779 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X780 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X781 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X782 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X783 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X784 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X785 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X786 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X787 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X788 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X789 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X790 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X791 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X792 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X793 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X794 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X795 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X796 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X797 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X798 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X799 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X800 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X801 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X802 tapered_buf_2/a_160_n140# tapered_buf_2/in tapered_buf_2/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X803 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X804 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X805 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X806 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X807 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X808 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X809 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X810 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X811 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X812 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X813 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X814 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X815 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X816 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X817 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X818 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X819 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X820 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X821 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X822 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X823 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X824 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X825 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X826 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X827 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X828 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X829 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X830 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X831 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X832 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X833 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X834 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X835 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X836 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X837 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X838 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X839 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X840 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X841 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X842 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X843 tapered_buf_2/a_580_0# tapered_buf_2/a_160_n140# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X844 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X845 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X846 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X847 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X848 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X849 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X850 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X851 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X852 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X853 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X854 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X855 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X856 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X857 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X858 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X859 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X860 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X861 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X862 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X863 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X864 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X865 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X866 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X867 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X868 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X869 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X870 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X871 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X872 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X873 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X874 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X875 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X876 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X877 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X878 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X879 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X880 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X881 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X882 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X883 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X884 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X885 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X886 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X887 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X888 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X889 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X890 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X891 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X892 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X893 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X894 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X895 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X896 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X897 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X898 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X899 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X900 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X901 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X902 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X903 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X904 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X905 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X906 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X907 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X908 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X909 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X910 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X911 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X912 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X913 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X914 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X915 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X916 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X917 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X918 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X919 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X920 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X921 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X922 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X923 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X924 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X925 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X926 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X927 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X928 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X929 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X930 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X931 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X932 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X933 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X934 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X935 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X936 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X937 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X938 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X939 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X940 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X941 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X942 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X943 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X944 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X945 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X946 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X947 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X948 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X949 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X950 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X951 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X952 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X953 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X954 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X955 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X956 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X957 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X958 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X959 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X960 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X961 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X962 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X963 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X964 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X965 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X966 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X967 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X968 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X969 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X970 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X971 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X972 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X973 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X974 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X975 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X976 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X977 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X978 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X979 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X980 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X981 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X982 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X983 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X984 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X985 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X986 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X987 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X988 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X989 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X990 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X991 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X992 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X993 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X994 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X995 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X996 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X997 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X998 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X999 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1000 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1001 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1002 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1003 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1004 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1005 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1006 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1007 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1008 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1009 gnd tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1010 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1011 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1012 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1013 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1014 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1015 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1016 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1017 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1018 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1019 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1020 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1021 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1022 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1023 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1024 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1025 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1026 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1027 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1028 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1029 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1030 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1031 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1032 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1034 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1035 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1036 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1037 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1038 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1039 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1040 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1041 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1042 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1043 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1044 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1045 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1046 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1047 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1048 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1049 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1050 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1051 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1052 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1053 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1055 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1056 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1057 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1058 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1059 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1060 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1061 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1062 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1063 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1064 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1065 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1066 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1067 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1068 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1069 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1070 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1071 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1072 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1073 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1074 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1075 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1076 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1077 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1078 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1079 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1080 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1081 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1082 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1083 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1084 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1085 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1086 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1087 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1088 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1089 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1090 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1091 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1092 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1093 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1094 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1095 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1096 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1097 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1098 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1099 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1100 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1101 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1102 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1103 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1104 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1105 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1106 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1107 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1108 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1109 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1110 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1111 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1112 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1113 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1114 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1115 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1116 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1117 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1118 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1119 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1120 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1121 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1122 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1123 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1124 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1125 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1126 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1127 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1128 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1129 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1130 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1131 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1132 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1133 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1134 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1135 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1136 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1137 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1138 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1139 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1140 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1141 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1142 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1143 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1144 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1145 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1146 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1147 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1148 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1149 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1150 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1151 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1152 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1153 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1154 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1155 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1156 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1157 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1158 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1159 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1160 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1161 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1162 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1163 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1164 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1165 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1166 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1167 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1168 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1169 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1170 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1171 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1172 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1173 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1174 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1175 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1176 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1177 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1178 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1179 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1180 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1181 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1182 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1183 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1184 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1185 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1186 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1187 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1188 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1189 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1190 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1191 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1192 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1193 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1194 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1195 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1196 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1197 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1198 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1199 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1200 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1201 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1202 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1203 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1204 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1205 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1206 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1207 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1208 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1209 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1210 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1211 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1212 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1213 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1214 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1215 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1216 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1217 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1218 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1219 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1220 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1221 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1222 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1223 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1224 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1225 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1226 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1227 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1228 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1229 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1230 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1231 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1232 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1233 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1234 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1235 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1236 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1237 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1238 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1239 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1240 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1241 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1242 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1243 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1244 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1245 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1246 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1247 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1248 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1249 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1250 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1251 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1252 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1253 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1254 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1255 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1256 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1257 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1258 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1259 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1260 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1261 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1262 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1263 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1264 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1265 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1266 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1267 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1268 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1269 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1270 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1271 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1272 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1273 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1274 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1275 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1276 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1277 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1278 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1279 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1280 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1281 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1282 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1283 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1284 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1285 gnd tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1286 tapered_buf_2/a_580_0# tapered_buf_2/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1287 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1288 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1289 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1290 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1291 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1292 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1293 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1294 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1295 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1296 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1297 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1298 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1299 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1300 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1301 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1302 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1303 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1304 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1305 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1306 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1307 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1308 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1309 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1310 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1311 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1312 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1313 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1314 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1315 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1316 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1317 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1318 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1319 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1320 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1321 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1322 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1323 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1324 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1326 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1327 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1328 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1329 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1330 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1331 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1332 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1333 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1334 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1335 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1336 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1337 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1338 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1339 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1340 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1341 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1342 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1343 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1344 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1345 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1346 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1347 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1348 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1349 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1350 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1351 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1352 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1353 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1354 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1355 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1356 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1357 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1358 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1359 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1360 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1361 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1362 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1363 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1364 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1365 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1366 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1367 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1368 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1369 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1370 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1371 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1372 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1373 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1374 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1375 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1376 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1377 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1378 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1379 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1380 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1381 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1382 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1383 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1384 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1385 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1386 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1387 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1388 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1389 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1390 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1391 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1392 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1393 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1394 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1395 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1396 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1397 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1398 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1399 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1400 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1401 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1402 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1403 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1404 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1405 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1406 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1407 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1408 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1409 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1410 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1411 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1412 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1413 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1414 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1415 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1416 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1417 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1418 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1419 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1420 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1421 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1422 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1423 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1424 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1425 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1426 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1427 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1428 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1429 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1430 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1431 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1432 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1433 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1434 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1435 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1436 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1437 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1438 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1439 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1440 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1441 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1442 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1443 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1444 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1445 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1446 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1447 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1448 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1449 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1450 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1451 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1452 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1453 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1454 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1455 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1456 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1457 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1458 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1459 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1460 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1461 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1462 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1463 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1464 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1465 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1466 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1467 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1468 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1469 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1470 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1471 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1472 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1473 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1474 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1475 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1476 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1477 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1478 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1479 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1480 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1481 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1482 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1483 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1484 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1485 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1486 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1487 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1488 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1489 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1490 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1491 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1492 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1493 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1494 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1495 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1496 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1497 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1498 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1499 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1500 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1501 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1502 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1503 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1504 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1505 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1506 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1507 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1508 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1509 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1510 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1511 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1512 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1513 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1514 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1515 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1516 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1517 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1518 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1519 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1520 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1521 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1522 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1523 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1524 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1525 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1526 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1527 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1528 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1529 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1530 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1531 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1532 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1533 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1534 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1535 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1536 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1537 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1538 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1539 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1540 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1541 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1542 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1543 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1544 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1545 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1546 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1547 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1548 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1549 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1550 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1551 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1552 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1553 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1554 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1555 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1556 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1557 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1558 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1559 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1560 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1561 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1562 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1563 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1564 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1565 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1566 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1567 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1568 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1569 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1570 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1571 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1572 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1573 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1574 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1575 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1576 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1577 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1578 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1579 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1580 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1581 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1582 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1583 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1584 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1585 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1586 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1587 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1588 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1589 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1590 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1591 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1592 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1593 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1594 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1595 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1596 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1597 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1598 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1599 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1600 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1601 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1602 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1603 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1604 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1605 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1606 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1607 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1608 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1610 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1611 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1612 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1613 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1614 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1615 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1616 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1617 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1618 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1619 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1620 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1621 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1622 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1623 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1624 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1625 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1626 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1627 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1628 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1629 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1630 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1631 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1632 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1633 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1634 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1635 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1636 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1637 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1638 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1639 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1640 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1641 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1642 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1643 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1644 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1645 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1646 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1647 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1648 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1649 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1650 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1651 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1652 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1653 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1654 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1655 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1656 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1657 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1658 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1659 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1660 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1661 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1662 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1663 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1664 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1665 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1666 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1667 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1668 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1669 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1670 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1671 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1672 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1673 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1674 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1675 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1676 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1677 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1678 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1679 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1680 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1681 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1682 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1683 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1684 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1685 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1686 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1687 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1688 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1689 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1690 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1691 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1692 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1693 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1694 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1695 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1696 gnd tapered_buf_2/a_210_n610# ro_complete_0/a5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1697 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1698 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1699 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1700 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1701 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1702 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1703 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1704 ro_complete_0/a5 tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1705 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1706 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1707 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1708 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1709 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1710 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1711 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1712 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1713 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1714 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1715 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1716 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1717 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1718 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1719 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1720 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1721 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1722 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1723 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1724 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1725 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1726 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1727 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1728 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1729 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1730 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1731 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1732 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1733 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1734 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1735 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1736 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1737 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1738 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1739 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1740 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1741 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1742 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1743 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1744 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1745 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1746 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1747 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1748 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1749 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1750 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1751 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1752 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1753 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1754 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1755 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1756 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1757 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1758 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1759 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1760 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1761 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1762 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1763 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1764 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1765 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1766 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1767 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1768 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1769 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1770 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1771 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1772 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1773 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1774 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1775 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1776 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1777 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1778 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1779 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1780 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1781 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1782 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1783 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1784 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1785 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1786 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1787 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1788 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1789 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1790 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1791 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1792 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1793 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1794 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1795 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1796 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1797 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1798 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1799 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1800 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1801 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1802 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1803 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1804 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1805 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1806 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1807 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1808 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1809 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1810 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1811 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1812 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1813 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1814 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1815 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1816 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1817 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1818 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1819 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1820 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1821 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1822 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1823 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1824 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1825 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1826 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1827 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1828 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1829 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1830 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1831 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1832 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1833 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1834 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1835 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1836 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1837 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1838 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1839 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1840 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1841 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1842 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1843 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1844 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1845 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1846 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1847 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1848 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1849 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1850 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1851 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1852 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1853 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1854 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1855 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1856 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1857 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1858 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1859 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1860 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1861 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1862 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1863 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1864 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1865 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1866 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1867 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1868 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1869 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1870 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1871 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1872 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1873 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1874 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1875 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1876 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1877 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1878 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1879 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1880 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1881 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1882 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1883 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1884 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1885 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1886 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1887 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1888 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1889 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1890 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1891 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1892 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1893 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1894 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1895 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1896 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1897 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1898 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1899 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1900 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1901 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1902 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1903 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1904 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1905 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1906 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1907 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1908 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1909 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1910 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1911 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1912 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1913 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1914 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1915 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1916 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1917 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1918 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1919 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1920 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1921 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1922 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1923 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1924 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1925 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1926 tapered_buf_3/a_160_230# tapered_buf_3/in tapered_buf_3/a_n10_230# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1927 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1928 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1929 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1930 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1931 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1932 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1933 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1934 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1935 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1936 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1937 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1938 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1939 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1940 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1941 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1942 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1943 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1944 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1945 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1946 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1947 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1948 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1949 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1950 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1951 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1952 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1953 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1954 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1955 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1956 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1957 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1958 tapered_buf_3/a_580_0# tapered_buf_3/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1959 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1960 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1961 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1962 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1963 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1964 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1965 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1966 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1967 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1968 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1969 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1970 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1971 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1972 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1973 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1974 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1975 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1976 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1977 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1978 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1979 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1980 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1981 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1982 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1983 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1984 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1985 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1986 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1987 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1988 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1989 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1990 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1991 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1992 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1993 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1994 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1995 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1996 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1997 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1998 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1999 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2000 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2001 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2002 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2003 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2004 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2005 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2006 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2007 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2008 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2009 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2010 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2011 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2012 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2013 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2014 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2015 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2016 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2017 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2018 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2019 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2020 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2021 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2022 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2023 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2024 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2025 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2026 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2027 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2028 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2029 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2030 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2031 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2032 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2033 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2034 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2035 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2036 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2037 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2038 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2039 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2040 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2041 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2042 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2043 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2044 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2045 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2046 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2047 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2048 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2049 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2050 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2051 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2052 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2053 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2054 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2055 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2056 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2057 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2058 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2059 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2060 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2061 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2062 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2063 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2064 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2065 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2066 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2067 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2068 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2069 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2070 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2071 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2072 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2073 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2074 gnd tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2075 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2076 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2077 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2078 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2079 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2080 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2081 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2082 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2083 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2084 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2085 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2086 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2087 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2088 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2089 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2090 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2091 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2092 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2093 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2094 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2095 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2096 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2097 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2098 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2099 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2100 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2101 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2102 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2103 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2104 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2105 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2106 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2107 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2108 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2109 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2110 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2111 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2112 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2113 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2114 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2115 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2116 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2117 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2118 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2119 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2120 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2121 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2122 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2123 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2124 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2125 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2126 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2127 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2128 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2129 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2130 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2131 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2132 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2133 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2134 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2135 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2136 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2137 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2138 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2139 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2140 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2141 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2142 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2143 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2144 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2145 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2146 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2147 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2148 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2149 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2150 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2151 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2152 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2153 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2154 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2155 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2156 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2157 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2158 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2159 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2160 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2161 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2162 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2163 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2164 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2165 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2166 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2167 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2168 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2169 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2170 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2171 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2172 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2173 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2174 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2175 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2176 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2177 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2178 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2179 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2180 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2181 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2182 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2183 gnd tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2184 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2185 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2186 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2187 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2188 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2189 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2190 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2191 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2192 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2193 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2194 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2195 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2196 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2197 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2198 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2199 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2200 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2201 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2202 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2203 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2204 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2205 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2206 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2207 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2208 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2209 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2210 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2211 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2212 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2213 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2214 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2215 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2216 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2217 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2218 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2219 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2220 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2221 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2222 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2223 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2224 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2225 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2226 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2227 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2228 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2229 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2230 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2231 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2232 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2233 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2234 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2235 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2236 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2237 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2238 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2239 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2240 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2241 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2242 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2243 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2244 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2245 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2246 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2247 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2248 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2249 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2250 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2251 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2252 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2253 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2254 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2255 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2256 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2257 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2258 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2259 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2260 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2261 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2262 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2263 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2264 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2265 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2266 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2267 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2268 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2269 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2270 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2271 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2272 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2273 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2274 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2275 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2276 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2277 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2278 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2279 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2280 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2281 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2282 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2283 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2284 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2285 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2286 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2287 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2288 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2289 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2290 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2291 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2292 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2293 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2294 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2295 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2296 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2297 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2298 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2299 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2300 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2301 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2302 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2303 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2304 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2305 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2306 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2307 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2308 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2309 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2310 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2311 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2312 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2313 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2314 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2315 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2316 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2317 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2318 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2319 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2320 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2321 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2322 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2323 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2324 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2325 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2326 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2327 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2328 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2329 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2330 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2331 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2332 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2333 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2334 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2335 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2336 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2337 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2338 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2339 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2340 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2341 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2342 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2343 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2344 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2345 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2346 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2347 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2348 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2349 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2350 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2351 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2352 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2353 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2354 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2355 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2356 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2357 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2358 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2359 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2360 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2361 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2362 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2363 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2364 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2365 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2366 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2367 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2368 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2369 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2370 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2371 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2372 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2373 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2374 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2375 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2376 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2377 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2378 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2379 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2380 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2381 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2382 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2383 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2384 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2385 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2386 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2387 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2388 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2389 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2390 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2391 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2392 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2393 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2394 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2395 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2396 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2397 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2398 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2399 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2400 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2401 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2402 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2403 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2404 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2405 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2406 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2407 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2408 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2409 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2410 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2411 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2412 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2413 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2414 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2415 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2416 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2417 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2418 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2419 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2420 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2421 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2422 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2423 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2424 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2425 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2426 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2427 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2428 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2429 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2430 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2431 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2432 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2433 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2434 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2435 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2436 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2437 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2438 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2439 tapered_buf_3/a_580_0# tapered_buf_3/a_160_n140# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2440 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2441 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2442 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2443 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2444 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2445 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2446 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2447 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2448 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2449 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2450 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2451 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2452 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2453 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2454 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2455 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2456 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2457 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2458 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2459 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2460 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2461 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2462 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2463 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2464 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2465 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2466 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2467 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2468 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2469 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2470 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2471 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2472 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2473 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2474 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2475 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2476 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2477 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2478 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2479 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2480 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2481 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2482 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2483 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2484 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2485 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2486 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2487 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2488 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2489 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2490 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2491 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2492 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2493 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2494 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2495 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2496 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2497 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2498 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2499 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2500 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2501 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2502 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2503 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2504 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2505 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2506 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2507 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2508 tapered_buf_3/a_160_n140# tapered_buf_3/in tapered_buf_3/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2509 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2510 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2511 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2512 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2513 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2514 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2515 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2516 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2517 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2518 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2519 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2520 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2521 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2522 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2523 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2524 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2525 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2526 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2527 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2528 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2529 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2530 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2531 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2532 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2533 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2534 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2535 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2536 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2537 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2538 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2539 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2540 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2541 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2542 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2543 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2544 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2545 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2546 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2547 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2548 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2549 tapered_buf_3/a_580_0# tapered_buf_3/a_160_n140# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2550 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2551 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2552 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2553 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2554 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2555 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2556 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2557 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2558 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2559 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2560 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2561 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2562 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2563 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2564 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2565 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2566 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2567 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2568 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2569 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2570 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2571 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2572 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2573 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2574 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2575 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2576 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2577 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2578 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2579 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2580 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2581 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2582 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2583 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2584 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2585 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2586 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2587 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2588 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2589 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2590 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2591 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2592 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2593 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2594 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2595 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2596 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2597 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2598 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2599 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2600 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2601 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2602 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2603 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2604 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2605 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2606 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2607 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2608 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2609 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2610 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2611 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2612 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2613 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2614 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2615 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2616 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2617 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2618 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2619 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2620 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2621 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2622 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2623 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2624 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2625 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2626 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2627 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2628 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2629 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2630 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2631 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2632 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2633 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2634 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2635 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2636 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2637 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2638 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2639 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2640 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2641 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2642 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2643 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2644 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2645 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2646 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2647 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2648 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2649 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2650 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2651 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2652 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2653 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2654 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2655 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2656 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2657 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2658 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2659 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2660 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2661 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2662 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2663 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2664 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2665 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2666 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2667 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2668 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2669 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2670 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2671 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2672 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2673 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2674 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2675 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2676 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2677 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2678 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2679 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2680 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2681 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2682 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2683 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2684 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2685 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2686 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2687 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2688 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2689 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2690 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2691 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2692 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2693 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2694 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2695 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2696 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2697 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2698 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2699 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2700 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2701 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2702 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2703 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2704 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2705 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2706 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2707 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2708 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2709 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2710 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2711 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2712 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2713 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2714 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2715 gnd tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2716 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2717 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2718 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2719 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2720 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2721 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2722 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2723 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2724 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2725 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2726 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2727 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2728 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2729 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2730 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2731 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2732 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2733 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2734 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2735 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2736 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2737 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2738 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2739 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2740 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2741 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2742 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2743 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2744 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2745 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2746 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2747 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2748 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2749 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2750 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2751 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2752 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2753 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2754 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2755 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2756 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2757 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2758 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2759 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2760 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2761 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2762 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2763 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2764 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2765 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2766 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2767 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2768 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2769 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2770 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2771 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2772 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2773 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2774 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2775 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2776 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2777 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2778 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2779 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2780 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2781 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2782 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2783 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2784 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2785 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2786 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2787 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2788 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2789 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2790 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2791 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2792 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2793 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2794 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2795 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2796 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2797 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2798 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2799 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2800 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2801 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2802 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2803 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2804 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2805 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2806 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2807 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2808 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2809 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2810 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2811 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2812 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2813 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2814 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2815 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2816 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2817 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2818 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2819 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2820 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2821 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2822 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2823 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2824 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2825 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2826 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2827 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2828 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2829 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2830 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2831 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2832 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2833 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2834 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2835 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2836 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2837 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2838 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2839 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2840 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2841 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2842 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2843 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2844 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2845 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2846 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2847 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2848 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2849 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2850 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2851 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2852 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2853 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2854 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2855 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2856 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2857 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2858 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2859 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2860 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2861 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2862 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2863 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2864 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2865 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2866 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2867 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2868 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2869 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2870 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2871 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2872 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2873 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2874 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2875 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2876 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2877 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2878 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2879 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2880 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2881 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2882 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2883 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2884 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2885 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2886 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2887 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2888 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2889 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2890 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2891 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2892 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2893 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2894 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2895 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2896 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2897 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2898 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2899 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2900 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2901 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2902 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2903 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2904 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2905 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2906 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2907 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2908 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2909 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2910 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2911 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2912 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2913 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2914 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2915 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2916 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2917 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2918 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2919 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2920 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2921 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2922 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2923 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2924 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2925 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2926 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2927 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2928 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2929 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2930 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2931 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2932 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2933 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2934 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2935 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2936 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2937 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2938 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2939 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2940 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2941 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2942 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2943 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2944 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2945 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2946 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2947 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2948 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2949 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2950 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2951 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2952 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2953 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2954 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2955 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2956 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2957 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2958 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2959 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2960 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2961 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2962 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2963 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2964 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2965 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2966 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2967 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2968 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2969 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2970 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2971 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2972 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2973 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2974 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2975 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2976 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2977 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2978 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2979 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2980 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2981 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2982 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2983 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2984 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2985 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2986 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2987 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2988 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2989 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2990 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2991 gnd tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2992 tapered_buf_3/a_580_0# tapered_buf_3/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2993 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2994 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2995 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2996 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2997 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2998 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2999 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3000 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3001 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3002 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3003 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3004 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3005 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3006 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3007 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3008 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3009 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3010 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3011 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3012 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3013 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3014 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3015 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3016 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3017 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3018 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3019 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3020 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3021 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3022 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3023 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3024 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3025 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3026 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3027 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3028 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3029 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3030 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3031 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3032 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3033 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3034 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3035 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3036 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3037 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3038 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3039 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3040 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3041 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3042 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3043 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3044 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3045 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3046 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3047 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3048 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3049 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3050 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3051 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3052 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3053 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3054 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3055 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3056 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3057 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3058 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3059 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3060 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3061 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3062 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3063 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3064 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3065 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3066 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3067 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3068 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3069 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3070 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3071 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3072 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3073 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3074 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3075 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3076 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3077 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3078 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3079 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3080 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3081 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3082 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3083 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3084 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3085 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3086 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3087 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3088 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3089 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3090 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3091 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3092 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3093 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3094 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3095 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3096 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3097 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3098 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3099 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3100 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3101 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3102 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3103 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3104 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3105 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3106 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3107 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3108 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3109 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3110 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3111 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3112 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3113 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3114 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3115 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3116 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3117 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3118 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3119 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3120 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3121 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3122 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3123 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3124 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3125 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3126 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3127 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3128 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3129 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3130 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3131 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3132 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3133 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3134 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3135 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3136 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3137 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3138 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3139 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3140 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3141 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3142 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3143 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3144 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3145 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3146 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3147 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3148 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3149 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3150 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3151 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3152 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3153 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3154 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3155 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3156 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3157 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3158 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3159 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3160 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3161 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3162 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3163 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3164 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3165 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3166 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3167 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3168 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3169 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3170 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3171 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3172 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3173 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3174 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3175 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3176 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3177 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3178 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3179 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3180 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3181 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3182 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3183 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3184 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3185 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3186 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3187 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3188 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3189 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3190 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3191 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3192 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3193 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3194 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3195 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3196 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3197 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3198 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3199 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3200 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3201 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3202 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3203 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3204 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3205 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3206 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3207 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3208 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3209 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3210 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3211 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3212 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3213 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3214 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3215 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3216 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3217 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3218 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3219 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3220 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3221 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3222 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3223 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3224 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3225 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3226 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3227 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3228 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3229 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3230 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3231 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3232 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3233 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3234 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3235 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3236 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3237 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3238 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3239 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3240 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3241 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3242 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3243 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3244 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3245 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3246 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3247 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3248 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3249 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3250 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3251 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3252 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3253 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3254 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3255 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3256 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3257 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3258 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3259 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3260 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3261 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3262 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3263 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3264 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3265 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3266 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3267 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3268 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3269 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3270 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3271 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3272 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3273 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3274 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3275 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3276 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3277 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3278 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3279 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3280 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3281 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3282 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3283 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3284 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3285 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3286 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3287 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3288 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3289 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3290 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3291 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3292 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3293 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3294 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3295 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3296 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3297 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3298 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3299 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3300 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3301 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3302 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3303 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3304 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3305 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3306 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3307 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3308 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3309 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3310 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3311 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3312 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3313 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3314 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3315 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3316 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3317 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3318 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3319 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3320 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3321 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3322 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3323 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3324 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3325 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3326 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3327 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3328 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3329 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3330 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3331 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3332 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3333 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3334 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3335 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3336 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3337 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3338 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3339 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3340 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3341 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3342 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3343 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3344 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3345 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3346 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3347 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3348 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3349 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3350 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3351 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3352 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3353 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3354 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3355 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3356 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3357 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3358 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3359 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3360 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3361 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3362 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3363 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3364 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3365 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3366 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3367 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3368 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3369 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3370 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3371 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3372 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3373 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3374 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3375 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3376 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3377 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3378 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3379 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3380 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3381 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3382 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3383 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3384 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3385 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3386 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3387 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3388 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3389 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3390 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3391 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3392 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3393 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3394 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3395 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3396 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3397 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3398 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3399 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3400 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3401 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3402 gnd tapered_buf_3/a_210_n610# ro_complete_0/a4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3403 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3404 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3405 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3406 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3407 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3408 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3409 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3410 ro_complete_0/a4 tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3411 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3412 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3413 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3414 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3415 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3416 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3417 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3418 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3419 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3420 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3421 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3422 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3423 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3424 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3425 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3426 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3427 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3428 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3429 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3430 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3431 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3432 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3433 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3434 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3435 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3436 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3437 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3438 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3439 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3440 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3441 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3442 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3443 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3444 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3445 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3446 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3447 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3448 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3449 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3450 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3451 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3452 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3453 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3454 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3455 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3456 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3457 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3458 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3459 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3460 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3461 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3462 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3463 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3464 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3465 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3466 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3467 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3468 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3469 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3470 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3471 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3472 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3473 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3474 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3475 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3476 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3477 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3478 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3479 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3480 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3481 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3482 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3483 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3484 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3485 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3486 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3487 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3488 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3489 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3490 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3491 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3492 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3493 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3494 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3495 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3496 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3497 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3498 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3499 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3500 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3501 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3502 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3503 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3504 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3505 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3506 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3507 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3508 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3509 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3510 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3511 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3512 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3513 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3514 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3515 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3516 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3517 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3518 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3519 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3520 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3521 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3522 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3523 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3524 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3525 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3526 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3527 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3528 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3529 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3530 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3531 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3532 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3533 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3534 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3535 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3536 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3537 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3538 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3539 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3540 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3541 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3542 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3543 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3544 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3545 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3546 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3547 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3548 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3549 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3550 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3551 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3552 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3553 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3554 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3555 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3556 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3557 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3558 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3559 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3560 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3561 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3562 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3563 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3564 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3565 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3566 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3567 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3568 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3569 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3570 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3571 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3572 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3573 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3574 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3575 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3576 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3577 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3578 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3579 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3580 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3581 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3582 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3583 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3584 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3585 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3586 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3587 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3588 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3589 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3590 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3591 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3592 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3593 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3594 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3595 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3596 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3597 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3598 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3599 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3600 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3601 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3602 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3603 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3604 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3605 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3606 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3607 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3608 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3609 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3610 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3611 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3612 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3613 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3614 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3615 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3616 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3617 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3618 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3619 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3620 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3621 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3622 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3623 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3624 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3625 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3626 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3627 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3628 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3629 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3630 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3631 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3632 tapered_buf_4/a_160_230# tapered_buf_4/in tapered_buf_4/a_n10_230# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3633 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3634 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3635 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3636 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3637 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3638 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3639 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3640 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3641 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3642 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3643 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3644 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3645 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3646 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3647 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3648 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3649 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3650 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3651 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3652 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3653 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3654 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3655 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3656 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3657 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3658 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3659 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3660 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3661 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3662 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3663 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3664 tapered_buf_4/a_580_0# tapered_buf_4/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3665 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3666 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3667 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3668 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3669 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3670 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3671 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3672 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3673 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3674 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3675 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3676 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3677 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3678 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3679 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3680 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3681 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3682 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3683 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3684 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3685 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3686 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3687 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3688 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3689 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3690 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3691 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3692 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3693 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3694 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3695 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3696 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3697 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3698 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3699 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3700 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3701 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3702 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3703 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3704 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3705 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3706 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3707 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3708 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3709 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3710 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3711 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3712 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3713 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3714 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3715 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3716 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3717 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3718 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3719 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3720 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3721 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3722 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3723 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3724 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3725 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3726 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3727 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3728 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3729 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3730 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3731 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3732 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3733 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3734 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3735 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3736 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3737 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3738 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3739 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3740 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3741 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3742 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3743 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3744 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3745 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3746 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3747 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3748 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3749 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3750 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3751 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3752 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3753 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3754 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3755 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3756 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3757 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3758 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3759 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3760 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3761 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3762 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3763 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3764 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3765 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3766 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3767 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3768 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3769 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3770 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3771 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3772 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3773 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3774 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3775 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3776 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3777 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3778 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3779 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3780 gnd tapered_buf_4/a_160_n140# tapered_buf_4/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3781 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3782 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3783 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3784 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3785 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3786 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3787 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3788 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3789 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3790 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3791 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3792 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3793 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3794 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3795 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3796 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3797 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3798 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3799 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3800 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3801 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3802 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3803 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3804 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3805 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3806 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3807 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3808 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3809 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3810 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3811 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3812 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3813 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3814 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3815 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3816 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3817 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3818 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3819 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3820 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3821 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3822 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3823 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3824 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3825 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3826 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3827 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3828 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3829 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3830 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3831 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3832 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3833 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3834 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3835 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3836 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3837 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3838 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3839 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3840 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3841 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3842 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3843 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3844 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3845 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3846 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3847 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3848 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3849 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3850 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3851 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3852 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3853 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3854 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3855 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3856 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3857 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3858 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3859 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3860 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3861 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3862 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3863 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3864 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3865 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3866 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3867 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3868 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3869 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3870 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3871 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3872 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3873 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3874 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3875 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3876 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3877 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3878 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3879 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3880 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3881 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3882 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3883 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3884 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3885 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3886 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3887 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3888 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3889 gnd tapered_buf_4/a_160_n140# tapered_buf_4/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3890 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3891 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3892 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3893 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3894 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3895 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3896 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3897 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3898 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3899 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3900 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3901 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3902 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3903 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3904 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3905 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3906 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3907 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3908 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3909 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3910 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3911 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3912 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3913 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3914 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3915 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3916 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3917 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3918 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3919 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3920 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3921 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3922 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3923 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3924 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3925 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3926 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3927 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3928 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3929 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3930 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3931 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3932 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3933 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3934 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3935 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3936 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3937 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3938 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3939 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3940 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3941 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3942 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3943 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3944 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3945 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3946 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3947 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3948 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3949 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3950 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3951 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3952 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3953 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3954 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3955 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3956 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3957 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3958 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3959 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3960 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3961 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3962 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3963 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3964 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3965 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3966 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3967 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3968 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3969 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3970 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3971 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3972 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3973 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3974 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3975 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3976 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3977 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3978 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3979 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3980 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3981 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3982 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3983 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3984 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3985 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3986 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3987 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3988 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3989 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3990 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3991 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3992 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3993 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3994 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3995 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3996 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3997 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3998 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3999 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4000 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4001 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4002 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4003 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4004 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4005 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4006 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4007 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4008 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4009 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4010 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4011 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4012 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4013 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4014 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4015 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4016 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4017 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4018 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4019 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4020 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4021 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4022 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4023 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4024 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4025 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4026 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4027 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4028 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4029 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4030 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4031 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4032 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4033 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4034 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4035 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4036 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4037 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4038 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4039 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4040 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4041 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4042 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4043 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4044 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4045 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4046 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4047 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4048 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4049 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4050 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4051 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4052 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4053 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4054 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4055 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4056 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4057 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4058 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4059 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4060 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4061 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4062 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4063 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4064 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4065 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4066 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4067 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4068 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4069 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4070 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4071 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4072 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4073 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4074 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4075 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4076 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4077 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4078 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4079 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4080 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4081 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4082 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4083 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4084 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4085 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4086 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4087 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4088 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4089 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4090 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4091 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4092 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4093 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4094 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4095 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4096 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4097 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4098 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4099 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4100 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4101 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4102 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4103 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4104 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4105 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4106 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4107 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4108 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4109 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4110 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4111 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4112 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4113 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4114 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4115 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4116 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4117 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4118 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4119 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4120 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4121 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4122 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4123 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4124 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4125 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4126 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4127 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4128 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4129 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4130 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4131 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4132 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4133 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4134 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4135 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4136 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4137 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4138 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4139 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4140 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4141 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4142 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4143 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4144 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4145 tapered_buf_4/a_580_0# tapered_buf_4/a_160_n140# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4146 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4147 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4148 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4149 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4150 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4151 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4152 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4153 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4154 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4155 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4156 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4157 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4158 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4159 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4160 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4161 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4162 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4163 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4164 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4165 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4166 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4167 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4168 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4169 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4170 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4171 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4172 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4173 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4174 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4175 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4176 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4177 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4178 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4179 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4180 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4181 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4182 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4183 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4184 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4185 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4186 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4187 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4188 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4189 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4190 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4191 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4192 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4193 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4194 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4195 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4196 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4197 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4198 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4199 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4200 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4201 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4202 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4203 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4204 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4205 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4206 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4207 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4208 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4209 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4210 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4211 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4212 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4213 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4214 tapered_buf_4/a_160_n140# tapered_buf_4/in tapered_buf_4/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4215 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4216 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4217 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4218 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4219 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4220 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4221 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4222 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4223 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4224 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4225 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4226 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4227 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4228 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4229 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4230 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4231 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4232 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4233 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4234 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4235 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4236 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4237 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4238 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4239 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4240 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4241 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4242 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4243 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4244 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4245 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4246 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4247 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4248 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4249 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4250 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4251 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4252 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4253 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4254 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4255 tapered_buf_4/a_580_0# tapered_buf_4/a_160_n140# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4256 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4257 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4258 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4259 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4260 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4261 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4262 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4263 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4264 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4265 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4266 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4267 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4268 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4269 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4270 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4271 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4272 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4273 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4274 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4275 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4276 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4277 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4278 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4279 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4280 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4281 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4282 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4283 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4284 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4285 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4286 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4287 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4288 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4289 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4290 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4291 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4292 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4293 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4294 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4295 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4296 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4297 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4298 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4299 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4300 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4301 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4302 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4303 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4304 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4305 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4306 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4307 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4308 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4309 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4310 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4311 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4312 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4313 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4314 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4315 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4316 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4317 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4318 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4319 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4320 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4321 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4322 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4323 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4324 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4325 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4326 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4327 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4328 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4329 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4330 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4331 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4332 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4333 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4334 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4335 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4336 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4337 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4338 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4339 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4340 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4341 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4342 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4343 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4344 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4345 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4346 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4347 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4348 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4349 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4350 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4351 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4352 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4353 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4354 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4355 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4356 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4357 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4358 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4359 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4360 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4361 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4362 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4363 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4364 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4365 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4366 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4367 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4368 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4369 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4370 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4371 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4372 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4373 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4374 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4375 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4376 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4377 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4378 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4379 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4380 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4381 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4382 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4383 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4384 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4385 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4386 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4387 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4388 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4389 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4390 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4391 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4392 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4393 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4394 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4395 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4396 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4397 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4398 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4399 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4400 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4401 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4402 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4403 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4404 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4405 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4406 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4407 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4408 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4409 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4410 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4411 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4412 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4413 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4414 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4415 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4416 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4417 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4418 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4419 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4420 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4421 gnd tapered_buf_4/a_160_n140# tapered_buf_4/a_580_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4422 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4423 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4424 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4425 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4426 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4427 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4428 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4429 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4430 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4431 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4432 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4433 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4434 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4435 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4436 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4437 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4438 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4439 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4440 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4441 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4442 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4443 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4444 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4445 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4446 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4447 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4448 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4449 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4450 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4451 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4452 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4453 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4454 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4455 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4456 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4457 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4458 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4459 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4460 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4461 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4462 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4463 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4464 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4465 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4466 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4467 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4468 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4469 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4470 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4471 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4472 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4473 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4474 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4475 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4476 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4477 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4478 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4479 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4480 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4481 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4482 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4483 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4484 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4485 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4486 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4487 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4488 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4489 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4490 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4491 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4492 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4493 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4494 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4495 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4496 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4497 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4498 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4499 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4500 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4501 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4502 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4503 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4504 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4505 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4506 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4507 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4508 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4509 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4510 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4511 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4512 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4513 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4514 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4515 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4516 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4517 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4518 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4519 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4520 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4521 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4522 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4523 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4524 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4525 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4526 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4527 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4528 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4529 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4530 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4531 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4532 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4533 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4534 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4535 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4536 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4537 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4538 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4539 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4540 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4541 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4542 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4543 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4544 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4545 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4546 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4547 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4548 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4549 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4550 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4551 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4552 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4553 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4554 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4555 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4556 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4557 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4558 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4559 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4560 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4561 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4562 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4563 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4564 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4565 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4566 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4567 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4568 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4569 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4570 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4571 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4572 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4573 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4574 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4575 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4576 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4577 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4578 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4579 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4580 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4581 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4582 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4583 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4584 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4585 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4586 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4587 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4588 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4589 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4590 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4591 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4592 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4593 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4594 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4595 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4596 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4597 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4598 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4599 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4600 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4601 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4602 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4603 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4604 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4605 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4606 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4607 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4608 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4609 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4610 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4611 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4612 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4613 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4614 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4615 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4616 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4617 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4618 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4619 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4620 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4621 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4622 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4623 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4624 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4625 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4626 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4627 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4628 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4629 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4630 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4631 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4632 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4633 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4634 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4635 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4636 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4637 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4638 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4639 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4640 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4641 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4642 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4643 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4644 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4645 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4646 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4647 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4648 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4649 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4650 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4651 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4652 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4653 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4654 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4655 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4656 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4657 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4658 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4659 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4660 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4661 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4662 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4663 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4664 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4665 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4666 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4667 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4668 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4669 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4670 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4671 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4672 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4673 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4674 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4675 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4676 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4677 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4678 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4679 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4680 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4681 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4682 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4683 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4684 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4685 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4686 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4687 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4688 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4689 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4690 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4691 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4692 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4693 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4694 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4695 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4696 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4697 gnd tapered_buf_4/a_160_n140# tapered_buf_4/a_580_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4698 tapered_buf_4/a_580_0# tapered_buf_4/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4699 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4700 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4701 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4702 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4703 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4704 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4705 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4706 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4707 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4708 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4709 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4710 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4711 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4712 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4713 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4714 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4715 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4716 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4717 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4718 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4719 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4720 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4721 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4722 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4723 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4724 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4725 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4726 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4727 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4728 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4729 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4730 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4731 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4732 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4733 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4734 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4735 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4736 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4737 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4738 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4739 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4740 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4741 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4742 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4743 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4744 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4745 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4746 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4747 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4748 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4749 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4750 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4751 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4752 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4753 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4754 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4755 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4756 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4757 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4758 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4759 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4760 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4761 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4762 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4763 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4764 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4765 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4766 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4767 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4768 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4769 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4770 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4771 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4772 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4773 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4774 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4775 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4776 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4777 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4778 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4779 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4780 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4781 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4782 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4783 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4784 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4785 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4786 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4787 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4788 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4789 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4790 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4791 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4792 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4793 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4794 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4795 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4796 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4797 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4798 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4799 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4800 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4801 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4802 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4803 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4804 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4805 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4806 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4807 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4808 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4809 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4810 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4811 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4812 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4813 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4814 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4815 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4816 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4817 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4818 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4819 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4820 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4821 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4822 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4823 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4824 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4825 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4826 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4827 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4828 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4829 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4830 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4831 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4832 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4833 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4834 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4835 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4836 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4837 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4838 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4839 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4840 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4841 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4842 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4843 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4844 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4845 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4846 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4847 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4848 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4849 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4850 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4851 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4852 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4853 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4854 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4855 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4856 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4857 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4858 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4859 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4860 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4861 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4862 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4863 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4864 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4865 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4866 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4867 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4868 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4869 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4870 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4871 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4872 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4873 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4874 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4875 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4876 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4877 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4878 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4879 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4880 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4881 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4882 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4883 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4884 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4885 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4886 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4887 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4888 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4889 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4890 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4891 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4892 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4893 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4894 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4895 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4896 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4897 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4898 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4899 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4900 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4901 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4902 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4903 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4904 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4905 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4906 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4907 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4908 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4909 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4910 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4911 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4912 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4913 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4914 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4915 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4916 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4917 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4918 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4919 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4920 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4921 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4922 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4923 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4924 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4925 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4926 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4927 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4928 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4929 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4930 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4931 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4932 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4933 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4934 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4935 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4936 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4937 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4938 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4939 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4940 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4941 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4942 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4943 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4944 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4945 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4946 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4947 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4948 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4949 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4950 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4951 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4952 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4953 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4954 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4955 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4956 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4957 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4958 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4959 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4960 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4961 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4962 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4963 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4964 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4965 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4966 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4967 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4968 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4969 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4970 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4971 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4972 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4973 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4974 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4975 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4976 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4977 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4978 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4979 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4980 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4981 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4982 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4983 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4984 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4985 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4986 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4987 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4988 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4989 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4990 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4991 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4992 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4993 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4994 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4995 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4996 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4997 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4998 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4999 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5000 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5001 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5002 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5003 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5004 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5005 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5006 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5007 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5008 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5009 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5010 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5011 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5012 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5013 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5014 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5015 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5016 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5017 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5018 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5019 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5020 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5021 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5022 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5023 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5024 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5025 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5026 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5027 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5028 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5029 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5030 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5031 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5032 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5033 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5034 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5035 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5036 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5037 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5038 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5039 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5040 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5041 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5042 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5043 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5044 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5045 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5046 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5047 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5048 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5049 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5050 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5051 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5052 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5053 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5054 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5055 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5056 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5057 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5058 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5059 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5060 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5061 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5062 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5063 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5064 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5065 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5066 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5067 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5068 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5069 tapered_buf_4/a_1650_0# tapered_buf_4/a_580_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5070 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5071 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5072 gnd tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5073 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5074 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5075 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5076 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5077 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5078 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5079 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5080 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5081 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5082 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5083 gnd tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5084 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5085 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5086 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5087 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5088 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5089 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5090 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5091 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5092 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5093 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5094 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5095 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5096 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5097 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5098 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5099 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5100 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5101 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5102 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5103 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5104 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5105 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5106 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5107 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5108 gnd tapered_buf_4/a_210_n610# ro_complete_0/a3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5109 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5110 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5111 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5112 gnd tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# tapered_buf_4/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5113 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd tapered_buf_4/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5114 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5115 tapered_buf_4/a_210_n610# tapered_buf_4/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5116 ro_complete_0/a3 tapered_buf_4/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5117 tapered_buf_4/a_4670_0# tapered_buf_4/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5118 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5119 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5120 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5121 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5122 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5123 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5124 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5125 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5126 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5127 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5128 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5129 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5130 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5131 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5132 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5133 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5134 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5135 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5136 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5137 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5138 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5139 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5140 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5141 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5142 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5143 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5144 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5145 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5146 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5147 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5148 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5149 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5150 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5151 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5152 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5153 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5154 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5155 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5156 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5157 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5158 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5159 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5160 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5161 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5162 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5163 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5164 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5165 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5166 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5167 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5168 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5169 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5170 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5171 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5172 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5173 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5174 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5175 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5176 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5177 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5178 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5179 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5180 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5181 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5182 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5183 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5184 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5185 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5186 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5187 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5188 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5189 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5190 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5191 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5192 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5193 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5194 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5195 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5196 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5197 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5198 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5199 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5200 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5201 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5202 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5203 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5204 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5205 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5206 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5207 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5208 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5209 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5210 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5211 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5212 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5213 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5214 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5215 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5216 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5217 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5218 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5219 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5220 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5221 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5222 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5223 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5224 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5225 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5226 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5227 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5228 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5229 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5230 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5231 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5232 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5233 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5234 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5235 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5236 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5237 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5238 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5239 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5240 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5241 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5242 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5243 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5244 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5245 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5246 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5247 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5248 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5249 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5250 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5251 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5252 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5253 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5254 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5255 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5256 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5257 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5258 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5259 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5260 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5261 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5262 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5263 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5264 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5265 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5266 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5267 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5268 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5269 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5270 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5271 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5272 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5273 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5274 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5275 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5276 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5277 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5278 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5279 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5280 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5281 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5282 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5283 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5284 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5285 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5286 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5287 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5288 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5289 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5290 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5291 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5292 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5293 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5294 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5295 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5296 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5297 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5298 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5299 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5300 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5301 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5302 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5303 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5304 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5305 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5306 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5307 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5308 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5309 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5310 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5311 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5312 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5313 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5314 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5315 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5316 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5317 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5318 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5319 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5320 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5321 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5322 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5323 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5324 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5325 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5326 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5327 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5328 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5329 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5330 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5331 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5332 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5333 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5334 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5335 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5336 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5337 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5338 tapered_buf_5/a_160_230# tapered_buf_5/in tapered_buf_5/a_n10_230# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5339 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5340 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5341 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5342 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5343 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5344 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5345 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5346 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5347 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5348 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5349 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5350 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5351 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5352 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5353 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5354 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5355 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5356 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5357 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5358 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5359 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5360 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5361 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5362 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5363 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5364 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5365 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5366 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5367 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5368 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5369 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5370 tapered_buf_5/a_580_0# tapered_buf_5/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5371 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5372 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5373 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5374 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5375 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5376 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5377 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5378 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5379 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5380 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5381 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5382 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5383 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5384 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5385 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5386 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5387 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5388 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5389 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5390 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5391 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5392 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5393 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5394 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5395 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5396 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5397 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5398 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5399 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5400 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5401 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5402 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5403 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5404 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5405 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5406 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5407 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5408 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5409 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5410 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5411 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5412 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5413 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5414 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5415 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5416 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5417 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5418 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5419 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5420 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5421 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5422 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5423 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5424 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5425 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5426 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5427 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5428 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5429 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5430 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5431 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5432 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5433 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5434 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5435 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5436 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5437 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5438 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5439 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5440 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5441 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5442 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5443 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5444 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5445 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5446 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5447 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5448 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5449 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5450 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5451 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5452 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5453 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5454 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5455 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5456 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5457 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5458 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5459 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5460 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5461 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5462 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5463 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5464 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5465 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5466 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5467 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5468 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5469 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5470 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5471 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5472 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5473 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5474 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5475 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5476 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5477 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5478 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5479 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5480 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5481 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5482 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5483 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5484 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5485 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5486 gnd tapered_buf_5/a_160_n140# tapered_buf_5/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5487 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5488 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5489 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5490 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5491 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5492 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5493 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5494 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5495 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5496 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5497 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5498 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5499 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5500 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5501 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5502 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5503 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5504 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5505 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5506 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5507 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5508 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5509 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5510 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5511 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5512 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5513 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5514 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5515 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5516 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5517 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5518 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5519 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5520 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5521 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5522 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5523 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5524 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5525 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5526 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5527 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5528 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5529 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5530 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5531 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5532 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5533 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5534 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5535 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5536 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5537 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5538 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5539 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5540 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5541 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5542 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5543 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5544 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5545 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5546 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5547 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5548 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5549 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5550 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5551 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5552 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5553 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5554 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5555 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5556 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5557 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5558 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5559 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5560 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5561 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5562 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5563 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5564 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5565 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5566 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5567 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5568 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5569 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5570 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5571 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5572 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5573 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5574 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5575 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5576 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5577 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5578 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5579 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5580 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5581 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5582 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5583 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5584 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5585 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5586 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5587 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5588 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5589 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5590 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5591 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5592 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5593 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5594 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5595 gnd tapered_buf_5/a_160_n140# tapered_buf_5/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5596 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5597 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5598 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5599 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5600 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5601 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5602 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5603 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5604 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5605 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5606 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5607 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5608 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5609 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5610 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5611 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5612 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5613 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5614 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5615 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5616 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5617 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5618 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5619 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5620 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5621 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5622 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5623 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5624 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5625 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5626 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5627 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5628 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5629 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5630 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5631 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5632 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5633 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5634 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5635 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5636 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5637 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5638 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5639 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5640 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5641 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5642 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5643 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5644 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5645 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5646 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5647 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5648 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5649 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5650 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5651 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5652 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5653 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5654 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5655 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5656 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5657 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5658 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5659 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5660 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5661 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5662 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5663 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5664 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5665 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5666 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5667 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5668 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5669 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5670 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5671 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5672 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5673 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5674 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5675 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5676 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5677 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5678 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5679 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5680 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5681 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5682 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5683 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5684 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5685 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5686 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5687 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5688 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5689 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5690 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5691 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5692 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5693 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5694 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5695 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5696 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5697 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5698 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5699 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5700 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5701 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5702 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5703 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5704 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5705 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5706 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5707 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5708 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5709 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5710 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5711 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5712 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5713 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5714 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5715 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5716 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5717 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5718 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5719 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5720 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5721 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5722 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5723 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5724 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5725 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5726 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5727 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5728 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5729 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5730 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5731 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5732 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5733 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5734 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5735 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5736 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5737 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5738 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5739 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5740 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5741 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5742 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5743 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5744 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5745 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5746 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5747 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5748 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5749 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5750 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5751 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5752 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5753 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5754 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5755 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5756 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5757 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5758 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5759 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5760 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5761 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5762 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5763 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5764 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5765 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5766 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5767 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5768 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5769 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5770 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5771 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5772 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5773 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5774 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5775 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5776 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5777 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5778 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5779 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5780 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5781 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5782 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5783 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5784 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5785 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5786 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5787 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5788 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5789 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5790 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5791 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5792 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5793 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5794 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5795 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5796 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5797 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5798 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5799 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5800 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5801 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5802 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5803 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5804 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5805 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5806 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5807 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5808 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5809 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5810 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5811 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5812 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5813 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5814 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5815 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5816 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5817 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5818 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5819 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5820 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5821 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5822 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5823 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5824 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5825 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5826 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5827 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5828 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5829 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5830 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5831 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5832 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5833 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5834 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5835 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5836 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5837 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5838 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5839 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5840 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5841 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5842 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5843 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5844 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5845 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5846 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5847 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5848 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5849 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5850 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5851 tapered_buf_5/a_580_0# tapered_buf_5/a_160_n140# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5852 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5853 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5854 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5855 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5856 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5857 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5858 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5859 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5860 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5861 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5862 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5863 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5864 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5865 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5866 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5867 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5868 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5869 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5870 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5871 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5872 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5873 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5874 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5875 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5876 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5877 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5878 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5879 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5880 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5881 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5882 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5883 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5884 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5885 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5886 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5887 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5888 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5889 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5890 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5891 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5892 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5893 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5894 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5895 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5896 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5897 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5898 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5899 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5900 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5901 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5902 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5903 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5904 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5905 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5906 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5907 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5908 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5909 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5910 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5911 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5912 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5913 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5914 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5915 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5916 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5917 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5918 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5919 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5920 tapered_buf_5/a_160_n140# tapered_buf_5/in tapered_buf_5/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5921 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5922 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5923 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5924 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5925 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5926 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5927 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5928 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5929 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5930 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5931 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5932 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5933 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5934 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5935 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5936 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5937 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5938 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5939 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5940 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5941 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5942 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5943 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5944 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5945 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5946 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5947 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5948 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5949 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5950 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5951 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5952 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5953 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5954 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5955 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5956 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5957 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5958 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5959 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5960 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5961 tapered_buf_5/a_580_0# tapered_buf_5/a_160_n140# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5962 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5963 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5964 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5965 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5966 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5967 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5968 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5969 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5970 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5971 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5972 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5973 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5974 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5975 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5976 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5977 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5978 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5979 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5980 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5981 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5982 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5983 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5984 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5985 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5986 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5987 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5988 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5989 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5990 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5991 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5992 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5993 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5994 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5995 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5996 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5997 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5998 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5999 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6000 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6001 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6002 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6003 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6004 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6005 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6006 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6007 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6008 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6009 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6010 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6011 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6012 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6013 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6014 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6015 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6016 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6017 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6018 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6019 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6020 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6021 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6022 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6023 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6024 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6025 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6026 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6027 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6028 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6029 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6030 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6031 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6032 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6033 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6034 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6035 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6036 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6037 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6038 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6039 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6040 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6041 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6042 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6043 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6044 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6045 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6046 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6047 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6048 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6049 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6050 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6051 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6052 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6053 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6054 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6055 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6056 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6057 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6058 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6059 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6060 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6061 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6062 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6063 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6064 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6065 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6066 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6067 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6068 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6069 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6070 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6071 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6072 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6073 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6074 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6075 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6076 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6077 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6078 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6079 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6080 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6081 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6082 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6083 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6084 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6085 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6086 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6087 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6088 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6089 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6090 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6091 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6092 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6093 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6094 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6095 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6096 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6097 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6098 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6099 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6100 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6101 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6102 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6103 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6104 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6105 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6106 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6107 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6108 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6109 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6110 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6111 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6112 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6113 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6114 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6115 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6116 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6117 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6118 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6119 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6120 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6121 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6122 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6123 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6124 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6125 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6126 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6127 gnd tapered_buf_5/a_160_n140# tapered_buf_5/a_580_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6128 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6129 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6130 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6131 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6132 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6133 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6134 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6135 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6136 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6137 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6138 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6139 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6140 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6141 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6142 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6143 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6144 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6145 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6146 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6147 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6148 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6149 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6150 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6151 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6152 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6153 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6154 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6155 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6156 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6157 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6158 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6159 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6160 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6161 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6162 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6163 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6164 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6165 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6166 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6167 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6168 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6169 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6170 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6171 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6172 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6173 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6174 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6175 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6176 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6177 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6178 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6179 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6180 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6181 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6182 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6183 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6184 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6185 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6186 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6187 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6188 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6189 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6190 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6191 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6192 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6193 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6194 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6195 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6196 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6197 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6198 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6199 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6200 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6201 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6202 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6203 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6204 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6205 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6206 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6207 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6208 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6209 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6210 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6211 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6212 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6213 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6214 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6215 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6216 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6217 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6218 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6219 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6220 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6221 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6222 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6223 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6224 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6225 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6226 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6227 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6228 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6229 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6230 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6231 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6232 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6233 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6234 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6235 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6236 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6237 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6238 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6239 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6240 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6241 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6242 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6243 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6244 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6245 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6246 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6247 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6248 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6249 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6250 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6251 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6252 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6253 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6254 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6255 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6256 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6257 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6258 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6259 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6260 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6261 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6262 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6263 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6264 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6265 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6266 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6267 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6268 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6269 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6270 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6271 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6272 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6273 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6274 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6275 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6276 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6277 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6278 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6279 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6280 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6281 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6282 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6283 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6284 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6285 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6286 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6287 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6288 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6289 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6290 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6291 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6292 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6293 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6294 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6295 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6296 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6297 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6298 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6299 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6300 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6301 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6302 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6303 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6304 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6305 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6306 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6307 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6308 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6309 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6310 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6311 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6312 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6313 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6314 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6315 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6316 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6317 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6318 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6319 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6320 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6321 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6322 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6323 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6324 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6325 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6326 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6327 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6328 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6329 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6330 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6331 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6332 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6333 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6334 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6335 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6336 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6337 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6338 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6339 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6340 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6341 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6342 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6343 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6344 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6345 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6346 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6347 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6348 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6349 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6350 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6351 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6352 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6353 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6354 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6355 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6356 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6357 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6358 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6359 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6360 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6361 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6362 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6363 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6364 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6365 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6366 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6367 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6368 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6369 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6370 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6371 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6372 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6373 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6374 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6375 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6376 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6377 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6378 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6379 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6380 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6381 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6382 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6383 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6384 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6385 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6386 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6387 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6388 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6389 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6390 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6391 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6392 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6393 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6394 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6395 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6396 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6397 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6398 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6399 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6400 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6401 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6402 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6403 gnd tapered_buf_5/a_160_n140# tapered_buf_5/a_580_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6404 tapered_buf_5/a_580_0# tapered_buf_5/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6405 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6406 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6407 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6408 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6409 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6410 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6411 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6412 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6413 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6414 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6415 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6416 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6417 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6418 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6419 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6420 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6421 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6422 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6423 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6424 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6425 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6426 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6427 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6428 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6429 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6430 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6431 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6432 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6433 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6434 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6435 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6436 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6437 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6438 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6439 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6440 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6441 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6442 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6443 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6444 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6445 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6446 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6447 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6448 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6449 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6450 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6451 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6452 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6453 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6454 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6455 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6456 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6457 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6458 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6459 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6460 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6461 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6462 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6463 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6464 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6465 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6466 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6467 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6468 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6469 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6470 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6471 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6472 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6473 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6474 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6475 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6476 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6477 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6478 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6479 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6480 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6481 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6482 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6483 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6484 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6485 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6486 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6487 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6488 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6489 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6490 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6491 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6492 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6493 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6494 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6495 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6496 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6497 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6498 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6499 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6500 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6501 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6502 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6503 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6504 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6505 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6506 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6507 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6508 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6509 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6510 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6511 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6512 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6513 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6514 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6515 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6516 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6517 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6518 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6519 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6520 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6521 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6522 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6523 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6524 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6525 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6526 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6527 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6528 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6529 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6530 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6531 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6532 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6533 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6534 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6535 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6536 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6537 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6538 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6539 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6540 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6541 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6542 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6543 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6544 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6545 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6546 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6547 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6548 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6549 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6550 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6551 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6552 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6553 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6554 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6555 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6556 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6557 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6558 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6559 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6560 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6561 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6562 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6563 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6564 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6565 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6566 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6567 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6568 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6569 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6570 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6571 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6572 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6573 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6574 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6575 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6576 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6577 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6578 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6579 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6580 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6581 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6582 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6583 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6584 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6585 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6586 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6587 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6588 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6589 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6590 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6591 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6592 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6593 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6594 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6595 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6596 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6597 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6598 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6599 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6600 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6601 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6602 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6603 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6604 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6605 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6606 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6607 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6608 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6609 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6610 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6611 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6612 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6613 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6614 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6615 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6616 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6617 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6618 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6619 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6620 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6621 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6622 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6623 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6624 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6625 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6626 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6627 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6628 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6629 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6630 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6631 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6632 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6633 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6634 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6635 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6636 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6637 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6638 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6639 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6640 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6641 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6642 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6643 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6644 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6645 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6646 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6647 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6648 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6649 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6650 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6651 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6652 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6653 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6654 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6655 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6656 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6657 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6658 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6659 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6660 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6661 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6662 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6663 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6664 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6665 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6666 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6667 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6668 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6669 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6670 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6671 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6672 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6673 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6674 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6675 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6676 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6677 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6678 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6679 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6680 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6681 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6682 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6683 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6684 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6685 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6686 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6687 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6688 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6689 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6690 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6691 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6692 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6693 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6694 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6695 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6696 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6697 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6698 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6699 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6700 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6701 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6702 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6703 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6704 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6705 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6706 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6707 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6708 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6709 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6710 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6711 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6712 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6713 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6714 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6715 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6716 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6717 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6718 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6719 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6720 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6721 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6722 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6723 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6724 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6725 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6726 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6727 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6728 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6729 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6730 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6731 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6732 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6733 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6734 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6735 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6736 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6737 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6738 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6739 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6740 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6741 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6742 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6743 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6744 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6745 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6746 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6747 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6748 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6749 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6750 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6751 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6752 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6753 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6754 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6755 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6756 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6757 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6758 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6759 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6760 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6761 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6762 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6763 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6764 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6765 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6766 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6767 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6768 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6769 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6770 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6771 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6772 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6773 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6774 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6775 tapered_buf_5/a_1650_0# tapered_buf_5/a_580_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6776 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6777 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6778 gnd tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6779 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6780 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6781 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6782 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6783 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6784 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6785 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6786 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6787 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6788 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6789 gnd tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6790 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6791 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6792 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6793 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6794 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6795 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6796 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6797 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6798 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6799 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6800 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6801 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6802 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6803 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6804 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6805 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6806 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6807 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6808 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6809 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6810 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6811 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6812 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6813 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6814 gnd tapered_buf_5/a_210_n610# ro_complete_0/a2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6815 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6816 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6817 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6818 gnd tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# tapered_buf_5/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6819 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd tapered_buf_5/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6820 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6821 tapered_buf_5/a_210_n610# tapered_buf_5/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6822 ro_complete_0/a2 tapered_buf_5/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6823 tapered_buf_5/a_4670_0# tapered_buf_5/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6824 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6825 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6826 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6827 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6828 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6829 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6830 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6831 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6832 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6833 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6834 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6835 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6836 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6837 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6838 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6839 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6840 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6841 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6842 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6843 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6844 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6845 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6846 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6847 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6848 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6849 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6850 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6851 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6852 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6853 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6854 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6855 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6856 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6857 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6858 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6859 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6860 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6861 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6862 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6863 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6864 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6865 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6866 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6867 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6868 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6869 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6870 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6871 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6872 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6873 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6874 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6875 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6876 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6877 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6878 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6879 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6880 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6881 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6882 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6883 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6884 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6885 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6886 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6887 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6888 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6889 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6890 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6891 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6892 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6893 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6894 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6895 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6896 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6897 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6898 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6899 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6900 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6901 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6902 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6903 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6904 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6905 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6906 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6907 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6908 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6909 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6910 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6911 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6912 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6913 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6914 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6915 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6916 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6917 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6918 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6919 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6920 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6921 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6922 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6923 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6924 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6925 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6926 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6927 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6928 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6929 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6930 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6931 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6932 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6933 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6934 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6935 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6936 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6937 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6938 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6939 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6940 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6941 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6942 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6943 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6944 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6945 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6946 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6947 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6948 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6949 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6950 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6951 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6952 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6953 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6954 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6955 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6956 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6957 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6958 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6959 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6960 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6961 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6962 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6963 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6964 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6965 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6966 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6967 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6968 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6969 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6970 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6971 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6972 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6973 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6974 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6975 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6976 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6977 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6978 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6979 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6980 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6981 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6982 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6983 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6984 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6985 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6986 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6987 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6988 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6989 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6990 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6991 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6992 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6993 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6994 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6995 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6996 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6997 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6998 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6999 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7000 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7001 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7002 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7003 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7004 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7005 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7006 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7007 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7008 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7009 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7010 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7011 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7012 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7013 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7014 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7015 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7016 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7017 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7018 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7019 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7020 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7021 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7022 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7023 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7024 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7025 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7026 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7027 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7028 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7029 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7030 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7031 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7032 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7033 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7034 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7035 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7036 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7037 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7038 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7039 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7040 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7041 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7042 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7043 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7044 tapered_buf_6/a_160_230# tapered_buf_6/in tapered_buf_6/a_n10_230# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7045 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7046 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7047 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7048 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7049 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7050 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7051 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7052 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7053 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7054 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7055 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7056 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7057 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7058 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7059 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7060 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7061 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7062 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7063 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7064 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7065 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7066 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7067 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7068 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7069 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7070 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7071 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7072 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7073 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7074 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7075 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7076 tapered_buf_6/a_580_0# tapered_buf_6/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7077 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7078 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7079 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7080 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7081 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7082 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7083 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7084 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7085 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7086 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7087 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7088 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7089 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7090 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7091 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7092 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7093 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7094 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7095 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7096 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7097 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7098 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7099 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7100 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7101 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7102 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7103 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7104 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7105 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7106 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7107 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7108 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7109 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7110 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7111 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7112 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7113 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7114 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7115 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7116 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7117 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7118 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7119 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7120 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7121 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7122 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7123 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7124 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7125 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7126 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7127 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7128 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7129 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7130 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7131 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7132 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7133 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7134 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7135 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7136 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7137 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7138 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7139 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7140 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7141 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7142 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7143 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7144 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7145 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7146 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7147 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7148 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7149 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7150 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7151 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7152 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7153 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7154 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7155 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7156 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7157 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7158 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7159 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7160 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7161 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7162 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7163 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7164 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7165 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7166 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7167 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7168 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7169 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7170 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7171 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7172 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7173 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7174 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7175 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7176 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7177 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7178 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7179 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7180 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7181 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7182 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7183 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7184 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7185 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7186 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7187 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7188 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7189 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7190 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7191 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7192 gnd tapered_buf_6/a_160_n140# tapered_buf_6/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7193 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7194 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7195 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7196 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7197 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7198 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7199 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7200 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7201 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7202 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7203 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7204 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7205 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7206 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7207 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7208 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7209 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7210 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7211 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7212 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7213 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7214 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7215 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7216 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7217 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7218 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7219 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7220 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7221 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7222 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7223 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7224 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7225 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7226 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7227 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7228 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7229 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7230 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7231 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7232 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7233 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7234 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7235 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7236 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7237 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7238 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7239 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7240 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7241 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7242 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7243 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7244 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7245 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7246 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7247 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7248 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7249 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7250 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7251 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7252 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7253 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7254 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7255 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7256 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7257 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7258 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7259 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7260 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7261 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7262 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7263 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7264 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7265 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7266 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7267 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7268 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7269 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7270 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7271 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7272 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7273 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7274 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7275 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7276 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7277 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7278 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7279 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7280 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7281 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7282 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7283 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7284 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7285 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7286 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7287 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7288 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7289 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7290 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7291 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7292 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7293 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7294 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7295 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7296 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7297 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7298 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7299 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7300 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7301 gnd tapered_buf_6/a_160_n140# tapered_buf_6/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7302 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7303 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7304 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7305 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7306 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7307 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7308 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7309 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7310 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7311 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7312 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7313 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7314 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7315 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7316 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7317 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7318 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7319 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7320 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7321 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7322 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7323 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7324 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7325 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7326 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7327 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7328 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7329 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7330 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7331 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7332 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7333 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7334 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7335 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7336 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7337 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7338 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7339 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7340 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7341 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7342 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7343 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7344 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7345 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7346 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7347 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7348 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7349 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7350 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7351 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7352 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7353 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7354 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7355 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7356 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7357 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7358 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7359 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7360 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7361 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7362 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7363 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7364 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7365 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7366 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7367 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7368 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7369 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7370 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7371 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7372 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7373 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7374 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7375 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7376 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7377 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7378 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7379 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7380 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7381 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7382 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7383 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7384 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7385 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7386 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7387 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7388 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7389 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7390 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7391 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7392 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7393 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7394 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7395 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7396 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7397 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7398 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7399 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7400 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7401 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7402 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7403 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7404 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7405 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7406 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7407 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7408 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7409 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7410 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7411 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7412 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7413 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7414 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7415 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7416 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7417 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7418 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7419 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7420 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7421 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7422 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7423 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7424 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7425 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7426 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7427 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7428 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7429 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7430 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7431 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7432 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7433 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7434 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7435 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7436 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7437 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7438 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7439 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7440 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7441 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7442 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7443 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7444 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7445 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7446 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7447 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7448 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7449 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7450 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7451 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7452 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7453 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7454 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7455 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7456 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7457 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7458 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7459 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7460 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7461 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7462 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7463 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7464 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7465 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7466 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7467 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7468 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7469 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7470 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7471 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7472 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7473 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7474 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7475 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7476 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7477 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7478 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7479 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7480 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7481 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7482 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7483 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7484 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7485 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7486 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7487 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7488 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7489 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7490 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7491 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7492 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7493 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7494 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7495 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7496 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7497 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7498 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7499 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7500 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7501 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7502 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7503 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7504 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7505 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7506 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7507 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7508 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7509 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7510 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7511 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7512 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7513 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7514 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7515 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7516 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7517 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7518 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7519 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7520 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7521 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7522 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7523 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7524 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7525 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7526 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7527 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7528 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7529 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7530 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7531 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7532 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7533 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7534 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7535 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7536 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7537 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7538 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7539 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7540 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7541 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7542 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7543 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7544 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7545 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7546 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7547 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7548 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7549 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7550 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7551 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7552 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7553 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7554 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7555 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7556 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7557 tapered_buf_6/a_580_0# tapered_buf_6/a_160_n140# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7558 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7559 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7560 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7561 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7562 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7563 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7564 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7565 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7566 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7567 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7568 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7569 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7570 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7571 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7572 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7573 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7574 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7575 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7576 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7577 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7578 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7579 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7580 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7581 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7582 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7583 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7584 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7585 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7586 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7587 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7588 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7589 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7590 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7591 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7592 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7593 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7594 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7595 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7596 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7597 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7598 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7599 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7600 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7601 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7602 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7603 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7604 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7605 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7606 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7607 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7608 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7609 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7610 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7611 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7612 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7613 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7614 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7615 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7616 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7617 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7618 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7619 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7620 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7621 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7622 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7623 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7624 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7625 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7626 tapered_buf_6/a_160_n140# tapered_buf_6/in tapered_buf_6/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7627 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7628 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7629 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7630 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7631 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7632 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7633 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7634 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7635 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7636 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7637 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7638 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7639 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7640 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7641 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7642 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7643 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7644 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7645 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7646 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7647 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7648 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7649 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7650 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7651 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7652 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7653 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7654 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7655 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7656 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7657 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7658 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7659 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7660 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7661 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7662 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7663 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7664 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7665 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7666 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7667 tapered_buf_6/a_580_0# tapered_buf_6/a_160_n140# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7668 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7669 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7670 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7671 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7672 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7673 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7674 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7675 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7676 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7677 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7678 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7679 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7680 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7681 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7682 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7683 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7684 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7685 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7686 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7687 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7688 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7689 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7690 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7691 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7692 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7693 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7694 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7695 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7696 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7697 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7698 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7699 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7700 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7701 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7702 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7703 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7704 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7705 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7706 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7707 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7708 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7709 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7710 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7711 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7712 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7713 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7714 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7715 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7716 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7717 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7718 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7719 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7720 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7721 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7722 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7723 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7724 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7725 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7726 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7727 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7728 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7729 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7730 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7731 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7732 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7733 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7734 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7735 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7736 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7737 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7738 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7739 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7740 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7741 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7742 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7743 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7744 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7745 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7746 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7747 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7748 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7749 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7750 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7751 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7752 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7753 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7754 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7755 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7756 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7757 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7758 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7759 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7760 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7761 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7762 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7763 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7764 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7765 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7766 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7767 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7768 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7769 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7770 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7771 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7772 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7773 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7774 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7775 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7776 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7777 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7778 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7779 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7780 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7781 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7782 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7783 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7784 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7785 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7786 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7787 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7788 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7789 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7790 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7791 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7792 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7793 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7794 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7795 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7796 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7797 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7798 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7799 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7800 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7801 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7802 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7803 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7804 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7805 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7806 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7807 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7808 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7809 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7810 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7811 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7812 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7813 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7814 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7815 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7816 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7817 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7818 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7819 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7820 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7821 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7822 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7823 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7824 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7825 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7826 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7827 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7828 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7829 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7830 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7831 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7832 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7833 gnd tapered_buf_6/a_160_n140# tapered_buf_6/a_580_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7834 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7835 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7836 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7837 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7838 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7839 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7840 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7841 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7842 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7843 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7844 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7845 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7846 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7847 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7848 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7849 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7850 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7851 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7852 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7853 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7854 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7855 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7856 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7857 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7858 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7859 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7860 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7861 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7862 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7863 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7864 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7865 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7866 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7867 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7868 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7869 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7870 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7871 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7872 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7873 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7874 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7875 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7876 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7877 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7878 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7879 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7880 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7881 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7882 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7883 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7884 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7885 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7886 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7887 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7888 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7889 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7890 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7891 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7892 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7893 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7894 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7895 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7896 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7897 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7898 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7899 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7900 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7901 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7902 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7903 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7904 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7905 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7906 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7907 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7908 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7909 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7910 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7911 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7912 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7913 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7914 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7915 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7916 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7917 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7918 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7919 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7920 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7921 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7922 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7923 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7924 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7925 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7926 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7927 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7928 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7929 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7930 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7931 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7932 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7933 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7934 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7935 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7936 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7937 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7938 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7939 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7940 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7941 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7942 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7943 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7944 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7945 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7946 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7947 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7948 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7949 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7950 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7951 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7952 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7953 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7954 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7955 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7956 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7957 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7958 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7959 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7960 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7961 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7962 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7963 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7964 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7965 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7966 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7967 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7968 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7969 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7970 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7971 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7972 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7973 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7974 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7975 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7976 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7977 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7978 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7979 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7980 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7981 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7982 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7983 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7984 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7985 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7986 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7987 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7988 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7989 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7990 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7991 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7992 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X7993 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7994 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7995 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7996 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7997 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7998 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7999 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8000 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8001 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8002 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8003 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8004 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8005 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8006 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8007 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8008 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8009 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8010 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8011 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8012 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8013 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8014 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8015 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8016 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8017 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8018 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8019 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8020 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8021 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8022 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8023 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8024 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8025 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8026 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8027 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8028 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8029 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8030 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8031 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8032 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8033 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8034 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8035 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8036 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8037 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8038 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8039 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8040 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8041 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8042 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8043 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8044 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8045 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8046 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8047 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8048 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8049 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8050 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8051 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8052 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8053 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8054 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8055 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8056 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8057 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8058 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8059 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8060 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8061 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8062 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8063 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8064 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8065 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8066 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8067 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8068 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8069 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8070 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8071 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8072 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8073 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8074 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8075 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8076 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8077 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8078 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8079 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8080 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8081 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8082 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8083 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8084 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8085 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8086 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8087 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8088 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8089 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8090 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8091 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8092 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8093 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8094 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8095 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8096 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8097 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8098 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8099 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8100 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8101 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8102 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8103 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8104 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8105 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8106 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8107 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8108 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8109 gnd tapered_buf_6/a_160_n140# tapered_buf_6/a_580_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8110 tapered_buf_6/a_580_0# tapered_buf_6/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8111 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8112 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8113 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8114 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8115 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8116 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8117 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8118 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8119 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8120 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8121 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8122 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8123 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8124 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8125 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8126 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8127 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8128 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8129 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8130 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8131 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8132 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8133 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8134 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8135 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8136 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8137 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8138 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8139 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8140 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8141 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8142 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8143 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8144 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8145 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8146 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8147 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8148 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8149 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8150 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8151 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8152 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8153 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8154 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8155 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8156 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8157 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8158 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8159 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8160 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8161 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8162 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8163 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8164 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8165 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8166 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8167 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8168 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8169 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8170 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8171 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8172 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8173 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8174 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8175 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8176 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8177 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8178 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8179 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8180 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8181 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8182 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8183 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8184 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8185 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8186 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8187 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8188 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8189 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8190 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8191 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8192 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8193 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8194 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8195 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8196 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8197 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8198 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8199 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8200 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8201 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8202 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8203 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8204 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8205 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8206 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8207 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8208 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8209 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8210 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8211 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8212 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8213 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8214 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8215 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8216 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8217 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8218 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8219 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8220 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8221 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8222 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8223 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8224 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8225 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8226 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8227 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8228 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8229 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8230 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8231 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8232 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8233 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8234 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8235 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8236 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8237 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8238 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8239 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8240 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8241 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8242 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8243 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8244 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8245 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8246 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8247 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8248 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8249 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8250 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8251 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8252 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8253 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8254 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8255 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8256 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8257 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8258 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8259 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8260 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8261 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8262 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8263 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8264 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8265 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8266 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8267 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8268 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8269 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8270 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8271 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8272 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8273 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8274 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8275 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8276 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8277 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8278 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8279 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8280 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8281 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8282 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8283 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8284 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8285 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8286 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8287 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8288 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8289 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8290 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8291 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8292 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8293 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8294 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8295 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8296 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8297 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8298 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8299 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8300 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8301 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8302 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8303 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8304 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8305 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8306 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8307 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8308 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8309 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8310 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8311 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8312 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8313 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8314 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8315 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8316 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8317 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8318 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8319 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8320 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8321 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8322 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8323 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8324 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8325 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8326 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8327 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8328 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8329 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8330 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8331 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8332 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8333 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8334 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8335 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8336 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8337 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8338 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8339 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8340 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8341 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8342 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8343 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8344 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8345 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8346 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8347 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8348 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8349 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8350 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8351 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8352 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8353 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8354 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8355 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8356 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8357 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8358 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8359 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8360 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8361 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8362 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8363 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8364 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8365 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8366 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8367 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8368 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8369 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8370 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8371 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8372 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8373 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8374 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8375 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8376 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8377 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8378 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8379 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8380 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8381 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8382 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8383 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8384 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8385 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8386 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8387 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8388 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8389 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8390 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8391 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8392 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8393 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8394 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8395 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8396 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8397 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8398 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8399 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8400 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8401 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8402 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8403 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8404 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8405 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8406 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8407 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8408 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8409 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8410 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8411 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8412 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8413 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8414 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8415 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8416 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8417 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8418 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8419 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8420 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8421 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8422 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8423 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8424 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8425 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8426 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8427 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8428 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8429 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8430 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8431 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8432 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8433 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8434 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8435 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8436 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8437 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8438 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8439 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8440 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8441 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8442 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8443 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8444 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8445 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8446 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8447 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8448 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8449 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8450 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8451 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8452 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8453 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8454 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8455 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8456 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8457 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8458 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8459 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8460 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8461 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8462 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8463 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8464 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8465 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8466 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8467 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8468 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8469 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8470 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8471 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8472 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8473 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8474 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8475 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8476 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8477 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8478 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8479 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8480 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8481 tapered_buf_6/a_1650_0# tapered_buf_6/a_580_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8482 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8483 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8484 gnd tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8485 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8486 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8487 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8488 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8489 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8490 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8491 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8492 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8493 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8494 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8495 gnd tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8496 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8497 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8498 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8499 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8500 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8501 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8502 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8503 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8504 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8505 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8506 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8507 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8508 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8509 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8510 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8511 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8512 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8513 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8514 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8515 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8516 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8517 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8518 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8519 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8520 gnd tapered_buf_6/a_210_n610# ro_complete_0/a1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8521 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8522 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8523 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8524 gnd tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# tapered_buf_6/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8525 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd tapered_buf_6/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8526 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8527 tapered_buf_6/a_210_n610# tapered_buf_6/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8528 ro_complete_0/a1 tapered_buf_6/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8529 tapered_buf_6/a_4670_0# tapered_buf_6/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8530 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8531 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8532 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8533 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8534 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8535 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8536 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8537 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8538 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8539 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8540 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8541 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8542 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8543 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8544 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8545 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8546 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8547 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8548 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8549 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8550 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8551 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8552 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8553 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8554 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8555 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8556 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8557 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8558 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8559 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8560 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8561 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8562 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8563 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8564 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8565 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8566 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8567 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8568 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8569 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8570 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8571 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8572 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8573 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8574 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8575 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8576 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8577 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8578 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8579 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8580 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8581 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8582 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8583 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8584 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8585 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8586 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8587 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8588 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8589 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8590 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8591 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8592 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8593 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8594 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8595 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8596 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8597 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8598 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8599 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8600 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8601 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8602 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8603 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8604 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8605 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8606 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8607 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8608 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8609 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8610 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8611 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8612 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8613 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8614 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8615 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8616 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8617 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8618 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8619 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8620 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8621 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8622 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8623 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8624 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8625 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8626 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8627 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8628 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8629 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8630 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8631 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8632 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8633 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8634 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8635 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8636 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8637 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8638 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8639 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8640 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8641 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8642 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8643 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8644 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8645 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8646 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8647 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8648 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8649 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8650 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8651 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8652 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8653 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8654 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8655 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8656 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8657 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8658 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8659 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8660 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8661 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8662 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8663 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8664 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8665 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8666 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8667 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8668 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8669 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8670 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8671 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8672 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8673 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8674 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8675 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8676 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8677 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8678 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8679 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8680 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8681 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8682 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8683 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8684 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8685 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8686 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8687 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8688 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8689 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8690 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8691 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8692 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8693 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8694 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8695 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8696 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8697 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8698 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8699 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8700 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8701 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8702 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8703 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8704 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8705 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8706 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8707 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8708 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8709 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8710 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8711 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8712 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8713 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8714 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8715 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8716 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8717 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8718 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8719 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8720 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8721 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8722 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8723 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8724 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8725 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8726 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8727 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8728 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8729 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8730 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8731 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8732 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8733 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8734 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8735 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8736 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8737 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8738 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8739 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8740 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8741 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8742 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8743 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8744 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8745 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8746 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8747 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8748 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8749 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8750 tapered_buf_7/a_160_230# tapered_buf_7/in tapered_buf_7/a_n10_230# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8751 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8752 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8753 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8754 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8755 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8756 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8757 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8758 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8759 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8760 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8761 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8762 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8763 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8764 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8765 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8766 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8767 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8768 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8769 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8770 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8771 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8772 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8773 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8774 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8775 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8776 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8777 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8778 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8779 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8780 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8781 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8782 tapered_buf_7/a_580_0# tapered_buf_7/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8783 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8784 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8785 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8786 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8787 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8788 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8789 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8790 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8791 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8792 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8793 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8794 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8795 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8796 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8797 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8798 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8799 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8800 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8801 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8802 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8803 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8804 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8805 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8806 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8807 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8808 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8809 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8810 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8811 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8812 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8813 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8814 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8815 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8816 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8817 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8818 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8819 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8820 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8821 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8822 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8823 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8824 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8825 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8826 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8827 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8828 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8829 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8830 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8831 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8832 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8833 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8834 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8835 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8836 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8837 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8838 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8839 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8840 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8841 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8842 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8843 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8844 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8845 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8846 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8847 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8848 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8849 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8850 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8851 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8852 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8853 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8854 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8855 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8856 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8857 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8858 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8859 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8860 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8861 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8862 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8863 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8864 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8865 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8866 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8867 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8868 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8869 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8870 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8871 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8872 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8873 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8874 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8875 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8876 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8877 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8878 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8879 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8880 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8881 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8882 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8883 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8884 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8885 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8886 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8887 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8888 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8889 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8890 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8891 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8892 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8893 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8894 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8895 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8896 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8897 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8898 gnd tapered_buf_7/a_160_n140# tapered_buf_7/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8899 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8900 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8901 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8902 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8903 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8904 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8905 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8906 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8907 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8908 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8909 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8910 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8911 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8912 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8913 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8914 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8915 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8916 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8917 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8918 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8919 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8920 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8921 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8922 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8923 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8924 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8925 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8926 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8927 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8928 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8929 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8930 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8931 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8932 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8933 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8934 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8935 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8936 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8937 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8938 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8939 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8940 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8941 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8942 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8943 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8944 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8945 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8946 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8947 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8948 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8949 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8950 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8951 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8952 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8953 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8954 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8955 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8956 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8957 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8958 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8959 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8960 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8961 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8962 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8963 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8964 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8965 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8966 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8967 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8968 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8969 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8970 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8971 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8972 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8973 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8974 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8975 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8976 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8977 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8978 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8979 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8980 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8981 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8982 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8983 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8984 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8985 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8986 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8987 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8988 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8989 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8990 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8991 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8992 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8993 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8994 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8995 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8996 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8997 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8998 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8999 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9000 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9001 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9002 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9003 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9004 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9005 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9006 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9007 gnd tapered_buf_7/a_160_n140# tapered_buf_7/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9008 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9009 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9010 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9011 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9012 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9013 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9014 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9015 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9016 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9017 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9018 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9019 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9020 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9021 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9022 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9023 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9024 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9025 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9026 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9027 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9028 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9029 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9030 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9031 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9032 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9033 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9034 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9035 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9036 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9037 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9038 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9039 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9040 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9041 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9042 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9043 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9044 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9045 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9046 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9047 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9048 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9049 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9050 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9051 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9052 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9053 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9054 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9055 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9056 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9057 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9058 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9059 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9060 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9061 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9062 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9063 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9064 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9065 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9066 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9067 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9068 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9069 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9070 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9071 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9072 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9073 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9074 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9075 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9076 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9077 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9078 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9079 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9080 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9081 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9082 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9083 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9084 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9085 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9086 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9087 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9088 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9089 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9090 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9091 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9092 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9093 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9094 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9095 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9096 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9097 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9098 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9099 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9100 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9101 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9102 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9103 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9104 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9105 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9106 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9107 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9108 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9109 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9110 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9111 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9112 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9113 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9114 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9115 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9116 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9117 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9118 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9119 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9120 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9121 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9122 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9123 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9124 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9125 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9126 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9127 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9128 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9129 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9130 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9131 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9132 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9133 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9134 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9135 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9136 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9137 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9138 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9139 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9140 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9141 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9142 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9143 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9144 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9145 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9146 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9147 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9148 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9149 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9150 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9151 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9152 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9153 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9154 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9155 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9156 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9157 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9158 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9159 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9160 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9161 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9162 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9163 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9164 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9165 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9166 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9167 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9168 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9169 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9170 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9171 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9172 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9173 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9174 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9175 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9176 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9177 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9178 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9179 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9180 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9181 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9182 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9183 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9184 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9185 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9186 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9187 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9188 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9189 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9190 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9191 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9192 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9193 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9194 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9195 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9196 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9197 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9198 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9199 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9200 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9201 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9202 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9203 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9204 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9205 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9206 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9207 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9208 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9209 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9210 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9211 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9212 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9213 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9214 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9215 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9216 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9217 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9218 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9219 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9220 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9221 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9222 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9223 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9224 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9225 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9226 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9227 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9228 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9229 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9230 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9231 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9232 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9233 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9234 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9235 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9236 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9237 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9238 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9239 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9240 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9241 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9242 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9243 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9244 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9245 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9246 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9247 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9248 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9249 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9250 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9251 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9252 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9253 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9254 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9255 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9256 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9257 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9258 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9259 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9260 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9261 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9262 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9263 tapered_buf_7/a_580_0# tapered_buf_7/a_160_n140# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9264 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9265 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9266 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9267 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9268 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9269 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9270 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9271 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9272 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9273 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9274 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9275 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9276 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9277 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9278 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9279 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9280 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9281 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9282 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9283 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9284 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9285 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9286 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9287 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9288 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9289 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9290 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9291 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9292 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9293 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9294 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9295 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9296 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9297 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9298 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9299 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9300 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9301 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9302 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9303 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9304 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9305 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9306 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9307 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9308 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9309 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9310 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9311 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9312 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9313 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9314 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9315 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9316 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9317 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9318 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9319 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9320 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9321 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9322 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9323 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9324 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9325 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9326 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9327 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9328 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9329 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9330 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9331 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9332 tapered_buf_7/a_160_n140# tapered_buf_7/in tapered_buf_7/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9333 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9334 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9335 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9336 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9337 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9338 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9339 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9340 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9341 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9342 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9343 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9344 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9345 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9346 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9347 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9348 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9349 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9350 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9351 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9352 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9353 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9354 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9355 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9356 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9357 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9358 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9359 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9360 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9361 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9362 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9363 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9364 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9365 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9366 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9367 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9368 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9369 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9370 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9371 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9372 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9373 tapered_buf_7/a_580_0# tapered_buf_7/a_160_n140# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9374 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9375 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9376 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9377 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9378 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9379 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9380 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9381 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9382 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9383 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9384 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9385 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9386 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9387 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9388 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9389 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9390 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9391 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9392 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9393 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9394 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9395 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9396 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9397 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9398 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9399 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9400 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9401 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9402 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9403 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9404 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9405 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9406 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9407 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9408 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9409 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9410 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9411 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9412 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9413 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9414 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9415 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9416 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9417 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9418 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9419 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9420 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9421 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9422 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9423 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9424 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9425 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9426 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9427 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9428 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9429 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9430 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9431 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9432 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9433 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9434 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9435 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9436 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9437 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9438 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9439 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9440 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9441 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9442 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9443 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9444 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9445 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9446 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9447 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9448 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9449 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9450 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9451 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9452 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9453 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9454 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9455 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9456 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9457 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9458 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9459 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9460 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9461 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9462 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9463 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9464 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9465 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9466 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9467 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9468 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9469 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9470 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9471 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9472 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9473 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9474 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9475 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9476 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9477 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9478 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9479 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9480 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9481 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9482 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9483 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9484 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9485 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9486 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9487 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9488 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9489 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9490 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9491 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9492 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9493 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9494 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9495 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9496 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9497 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9498 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9499 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9500 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9501 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9502 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9503 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9504 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9505 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9506 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9507 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9508 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9509 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9510 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9511 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9512 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9513 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9514 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9515 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9516 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9517 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9518 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9519 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9520 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9521 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9522 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9523 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9524 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9525 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9526 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9527 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9528 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9529 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9530 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9531 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9532 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9533 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9534 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9535 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9536 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9537 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9538 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9539 gnd tapered_buf_7/a_160_n140# tapered_buf_7/a_580_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9540 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9541 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9542 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9543 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9544 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9545 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9546 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9547 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9548 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9549 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9550 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9551 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9552 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9553 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9554 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9555 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9556 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9557 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9558 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9559 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9560 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9561 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9562 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9563 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9564 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9565 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9566 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9567 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9568 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9569 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9570 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9571 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9572 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9573 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9574 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9575 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9576 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9577 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9578 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9579 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9580 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9581 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9582 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9583 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9584 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9585 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9586 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9587 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9588 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9589 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9590 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9591 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9592 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9593 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9594 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9595 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9596 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9597 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9598 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9599 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9600 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9601 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9602 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9603 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9604 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9605 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9606 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9607 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9608 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9609 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9610 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9611 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9612 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9613 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9614 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9615 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9616 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9617 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9618 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9619 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9620 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9621 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9622 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9623 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9624 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9625 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9626 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9627 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9628 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9629 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9630 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9631 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9632 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9633 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9634 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9635 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9636 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9637 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9638 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9639 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9640 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9641 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9642 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9643 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9644 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9645 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9646 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9647 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9648 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9649 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9650 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9651 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9652 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9653 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9654 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9655 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9656 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9657 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9658 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9659 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9660 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9661 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9662 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9663 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9664 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9665 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9666 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9667 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9668 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9669 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9670 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9671 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9672 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9673 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9674 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9675 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9676 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9677 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9678 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9679 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9680 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9681 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9682 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9683 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9684 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9685 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9686 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9687 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9688 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9689 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9690 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9691 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9692 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9693 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9694 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9695 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9696 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9697 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9698 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9699 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9700 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9701 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9702 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9703 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9704 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9705 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9706 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9707 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9708 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9709 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9710 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9711 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9712 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9713 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9714 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9715 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9716 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9717 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9718 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9719 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9720 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9721 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9722 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9723 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9724 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9725 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9726 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9727 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9728 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9729 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9730 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9731 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9732 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9733 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9734 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9735 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9736 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9737 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9738 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9739 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9740 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9741 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9742 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9743 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9744 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9745 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9746 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9747 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9748 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9749 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9750 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9751 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9752 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9753 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9754 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9755 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9756 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9757 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9758 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9759 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9760 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9761 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9762 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9763 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9764 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9765 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9766 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9767 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9768 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9769 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9770 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9771 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9772 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9773 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9774 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9775 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9776 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9777 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9778 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9779 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9780 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9781 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9782 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9783 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9784 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9785 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9786 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9787 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9788 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9789 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9790 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9791 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9792 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9793 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9794 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9795 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9796 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9797 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9798 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9799 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9800 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9801 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9802 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9803 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9804 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9805 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9806 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9807 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9808 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9809 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9810 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9811 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9812 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9813 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9814 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9815 gnd tapered_buf_7/a_160_n140# tapered_buf_7/a_580_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9816 tapered_buf_7/a_580_0# tapered_buf_7/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9817 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9818 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9819 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9820 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9821 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9822 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9823 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9824 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9825 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9826 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9827 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9828 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9829 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9830 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9831 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9832 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9833 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9834 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9835 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9836 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9837 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9838 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9839 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9840 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9841 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9842 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9843 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9844 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9845 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9846 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9847 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9848 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9849 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9850 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9851 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9852 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9853 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9854 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9855 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9856 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9857 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9858 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9859 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9860 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9861 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9862 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9863 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9864 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9865 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9866 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9867 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9868 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9869 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9870 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9871 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9872 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9873 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9874 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9875 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9876 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9877 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9878 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9879 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9880 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9881 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9882 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9883 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9884 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9885 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9886 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9887 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9888 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9889 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9890 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9891 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9892 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9893 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9894 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9895 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9896 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9897 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9898 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9899 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9900 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9901 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9902 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9903 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9904 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9905 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9906 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9907 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9908 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9909 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9910 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9911 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9912 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9913 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9914 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9915 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9916 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9917 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9918 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9919 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9920 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9921 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9922 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9923 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9924 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9925 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9926 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9927 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9928 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9929 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9930 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9931 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9932 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9933 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9934 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9935 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9936 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9937 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9938 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9939 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9940 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9941 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9942 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9943 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9944 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9945 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9946 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9947 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9948 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9949 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9950 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9951 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9952 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9953 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9954 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9955 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9956 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9957 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9958 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9959 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9960 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9961 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9962 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9963 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9964 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9965 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9966 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9967 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9968 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9969 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9970 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9971 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9972 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9973 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9974 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9975 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9976 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9977 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9978 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9979 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9980 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9981 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9982 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9983 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9984 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9985 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9986 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9987 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9988 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9989 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9990 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9991 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9992 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9993 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9994 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9995 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9996 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9997 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9998 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9999 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10000 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10001 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10002 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10003 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10004 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10005 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10006 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10007 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10008 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10009 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10010 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10011 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10012 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10013 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10014 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10015 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10016 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10017 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10018 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10019 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10020 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10021 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10022 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10023 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10024 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10025 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10026 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10027 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10028 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10029 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10030 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10031 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10032 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10033 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10034 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10035 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10036 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10037 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10038 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10039 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10040 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10041 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10042 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10043 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10044 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10045 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10046 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10047 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10048 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10049 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10050 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10051 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10052 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10053 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10054 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10055 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10056 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10057 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10058 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10059 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10060 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10061 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10062 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10063 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10064 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10065 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10066 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10067 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10068 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10069 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10070 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10071 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10072 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10073 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10074 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10075 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10076 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10077 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10078 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10079 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10080 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10081 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10082 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10083 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10084 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10085 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10086 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10087 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10088 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10089 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10090 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10091 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10092 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10093 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10094 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10095 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10096 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10097 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10098 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10099 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10100 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10101 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10102 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10103 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10104 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10105 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10106 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10107 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10108 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10109 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10110 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10111 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10112 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10113 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10114 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10115 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10116 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10117 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10118 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10119 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10120 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10121 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10122 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10123 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10124 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10125 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10126 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10127 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10128 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10129 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10130 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10131 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10132 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10133 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10134 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10135 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10136 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10137 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10138 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10139 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10140 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10141 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10142 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10143 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10144 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10145 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10146 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10147 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10148 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10149 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10150 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10151 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10152 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10153 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10154 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10155 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10156 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10157 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10158 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10159 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10160 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10161 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10162 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10163 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10164 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10165 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10166 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10167 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10168 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10169 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10170 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10171 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10172 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10173 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10174 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10175 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10176 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10177 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10178 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10179 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10180 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10181 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10182 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10183 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10184 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10185 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10186 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10187 tapered_buf_7/a_1650_0# tapered_buf_7/a_580_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10188 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10189 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10190 gnd tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10191 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10192 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10193 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10194 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10195 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10196 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10197 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10198 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10199 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10200 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10201 gnd tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10202 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10203 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10204 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10205 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10206 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10207 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10208 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10209 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10210 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10211 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10212 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10213 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10214 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10215 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10216 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10217 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10218 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10219 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10220 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10221 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10222 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10223 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10224 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10225 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10226 gnd tapered_buf_7/a_210_n610# ro_complete_0/a0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10227 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10228 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10229 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10230 gnd tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# tapered_buf_7/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10231 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd tapered_buf_7/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10232 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10233 tapered_buf_7/a_210_n610# tapered_buf_7/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10234 ro_complete_0/a0 tapered_buf_7/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10235 tapered_buf_7/a_4670_0# tapered_buf_7/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10236 ro_complete_0/cbank_0/v tapered_buf_0/out tapered_buf_0/out sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=1e+06u l=180000u
X10237 tapered_buf_1/in tapered_buf_0/out tapered_buf_0/out sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=1e+06u l=180000u
X10238 ro_complete_0/cbank_1/v ro_complete_0/cbank_0/v ro_complete_0/ro_var_extend_0/vdd ro_complete_0/ro_var_extend_0/vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X10239 tapered_buf_1/in ro_complete_0/cbank_1/v ro_complete_0/ro_var_extend_0/vdd ro_complete_0/ro_var_extend_0/vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X10240 ro_complete_0/cbank_0/v tapered_buf_1/in ro_complete_0/ro_var_extend_0/vdd ro_complete_0/ro_var_extend_0/vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X10241 ro_complete_0/cbank_1/v tapered_buf_0/out tapered_buf_0/out sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=1e+06u l=180000u
X10242 ro_complete_0/cbank_1/v ro_complete_0/cbank_0/v gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X10243 ro_complete_0/cbank_0/v tapered_buf_1/in gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X10244 tapered_buf_1/in ro_complete_0/cbank_1/v gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X10245 gnd ro_complete_0/a0 ro_complete_0/cbank_0/switch_0/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10246 gnd ro_complete_0/a1 ro_complete_0/cbank_0/switch_1/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10247 gnd ro_complete_0/a3 ro_complete_0/cbank_0/switch_3/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10248 gnd ro_complete_0/a2 ro_complete_0/cbank_0/switch_2/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10249 gnd ro_complete_0/a4 ro_complete_0/cbank_0/switch_4/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10250 gnd ro_complete_0/a5 ro_complete_0/cbank_0/switch_5/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10251 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_3/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10252 ro_complete_0/cbank_0/v gnd sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5.2e+06u
X10253 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_5/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10254 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_4/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10255 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_0/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10256 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_1/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10257 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_2/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10258 gnd ro_complete_0/a0 ro_complete_0/cbank_1/switch_0/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10259 gnd ro_complete_0/a1 ro_complete_0/cbank_1/switch_1/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10260 gnd ro_complete_0/a3 ro_complete_0/cbank_1/switch_3/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10261 gnd ro_complete_0/a2 ro_complete_0/cbank_1/switch_2/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10262 gnd ro_complete_0/a4 ro_complete_0/cbank_1/switch_4/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10263 gnd ro_complete_0/a5 ro_complete_0/cbank_1/switch_5/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10264 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_3/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10265 ro_complete_0/cbank_1/v gnd sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5.2e+06u
X10266 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_5/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10267 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_4/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10268 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_0/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10269 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_1/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10270 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_2/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10271 gnd ro_complete_0/a0 ro_complete_0/cbank_2/switch_0/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10272 gnd ro_complete_0/a1 ro_complete_0/cbank_2/switch_1/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10273 gnd ro_complete_0/a3 ro_complete_0/cbank_2/switch_3/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10274 gnd ro_complete_0/a2 ro_complete_0/cbank_2/switch_2/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10275 gnd ro_complete_0/a4 ro_complete_0/cbank_2/switch_4/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10276 gnd ro_complete_0/a5 ro_complete_0/cbank_2/switch_5/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X10277 tapered_buf_1/in ro_complete_0/cbank_2/switch_3/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10278 tapered_buf_1/in gnd sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5.2e+06u
X10279 tapered_buf_1/in ro_complete_0/cbank_2/switch_5/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10280 tapered_buf_1/in ro_complete_0/cbank_2/switch_4/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10281 tapered_buf_1/in ro_complete_0/cbank_2/switch_0/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10282 tapered_buf_1/in ro_complete_0/cbank_2/switch_1/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10283 tapered_buf_1/in ro_complete_0/cbank_2/switch_2/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X10284 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10285 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10286 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10287 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10288 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10289 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10290 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10291 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10292 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10293 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10294 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10295 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10296 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10297 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10298 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10299 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10300 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10301 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10302 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10303 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10304 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10305 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10306 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10307 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10308 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10309 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10310 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10311 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10312 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10313 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10314 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10315 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10316 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10317 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10318 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10319 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10320 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10321 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10322 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10323 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10324 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10325 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10326 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10327 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10328 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10329 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10330 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10331 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10332 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10333 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10334 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10335 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10336 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10337 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10338 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10339 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10340 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10341 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10342 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10343 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10344 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10345 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10346 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10347 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10348 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10349 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10350 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10351 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10352 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10353 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10354 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10355 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10356 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10357 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10358 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10359 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10360 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10361 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10362 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10363 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10364 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10365 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10366 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10367 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10368 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10369 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10370 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10371 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10372 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10373 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10374 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10375 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10376 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10377 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10378 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10379 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10380 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10381 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10382 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10383 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10384 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10385 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10386 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10387 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10388 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10389 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10390 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10391 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10392 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10393 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10394 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10395 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10396 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10397 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10398 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10399 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10400 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10401 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10402 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10403 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10404 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10405 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10406 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10407 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10408 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10409 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10410 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10411 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10412 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10413 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10414 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10415 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10416 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10417 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10418 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10419 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10420 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10421 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10422 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10423 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10424 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10425 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10426 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10427 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10428 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10429 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10430 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10431 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10432 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10433 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10434 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10435 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10436 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10437 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10438 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10439 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10440 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10441 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10442 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10443 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10444 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10445 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10446 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10447 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10448 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10449 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10450 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10451 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10452 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10453 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10454 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10455 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10456 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10457 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10458 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10459 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10460 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10461 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10462 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10463 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10464 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10465 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10466 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10467 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10468 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10469 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10470 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10471 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10472 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10473 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10474 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10475 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10476 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10477 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10478 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10479 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10480 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10481 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10482 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10483 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10484 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10485 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10486 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10487 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10488 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10489 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10490 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10491 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10492 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10493 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10494 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10495 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10496 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10497 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10498 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10499 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10500 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10501 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10502 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10503 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10504 tapered_buf_1/a_160_230# tapered_buf_1/in tapered_buf_1/a_n10_230# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10505 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10506 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10507 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10508 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10509 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10510 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10511 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10512 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10513 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10514 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10515 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10516 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10517 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10518 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10519 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10520 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10521 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10522 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10523 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10524 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10525 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10526 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10527 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10528 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10529 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10530 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10531 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10532 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10533 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10534 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10535 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10536 tapered_buf_1/a_580_0# tapered_buf_1/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10537 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10538 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10539 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10540 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10541 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10542 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10543 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10544 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10545 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10546 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10547 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10548 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10549 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10550 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10551 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10552 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10553 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10554 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10555 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10556 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10557 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10558 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10559 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10560 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10561 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10562 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10563 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10564 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10565 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10566 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10567 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10568 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10569 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10570 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10571 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10572 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10573 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10574 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10575 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10576 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10577 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10578 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10579 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10580 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10581 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10582 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10583 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10584 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10585 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10586 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10587 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10588 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10589 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10590 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10591 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10592 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10593 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10594 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10595 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10596 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10597 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10598 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10599 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10600 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10601 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10602 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10603 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10604 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10605 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10606 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10607 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10608 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10609 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10610 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10611 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10612 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10613 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10614 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10615 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10616 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10617 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10618 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10619 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10620 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10621 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10622 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10623 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10624 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10625 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10626 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10627 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10628 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10629 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10630 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10631 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10632 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10633 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10634 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10635 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10636 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10637 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10638 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10639 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10640 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10641 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10642 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10643 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10644 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10645 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10646 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10647 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10648 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10649 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10650 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10651 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10652 gnd tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10653 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10654 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10655 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10656 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10657 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10658 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10659 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10660 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10661 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10662 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10663 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10664 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10665 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10666 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10667 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10668 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10669 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10670 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10671 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10672 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10673 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10674 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10675 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10676 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10677 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10678 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10679 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10680 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10681 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10682 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10683 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10684 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10685 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10686 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10687 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10688 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10689 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10690 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10691 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10692 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10693 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10694 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10695 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10696 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10697 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10698 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10699 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10700 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10701 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10702 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10703 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10704 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10705 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10706 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10707 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10708 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10709 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10710 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10711 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10712 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10713 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10714 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10715 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10716 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10717 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10718 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10719 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10720 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10721 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10722 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10723 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10724 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10725 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10726 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10727 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10728 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10729 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10730 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10731 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10732 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10733 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10734 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10735 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10736 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10737 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10738 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10739 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10740 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10741 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10742 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10743 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10744 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10745 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10746 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10747 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10748 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10749 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10750 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10751 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10752 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10753 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10754 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10755 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10756 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10757 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10758 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10759 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10760 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10761 gnd tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10762 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10763 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10764 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10765 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10766 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10767 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10768 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10769 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10770 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10771 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10772 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10773 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10774 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10775 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10776 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10777 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10778 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10779 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10780 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10781 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10782 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10783 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10784 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10785 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10786 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10787 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10788 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10789 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10790 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10791 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10792 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10793 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10794 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10795 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10796 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10797 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10798 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10799 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10800 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10801 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10802 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10803 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10804 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10805 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10806 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10807 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10808 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10809 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10810 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10811 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10812 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10813 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10814 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10815 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10816 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10817 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10818 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10819 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10820 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10821 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10822 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10823 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10824 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10825 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10826 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10827 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10828 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10829 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10830 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10831 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10832 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10833 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10834 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10835 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10836 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10837 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10838 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10839 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10840 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10841 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10842 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10843 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10844 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10845 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10846 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10847 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10848 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10849 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10850 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10851 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10852 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10853 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10854 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10855 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10856 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10857 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10858 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10859 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10860 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10861 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10862 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10863 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10864 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10865 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10866 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10867 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10868 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10869 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10870 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10871 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10872 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10873 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10874 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10875 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10876 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10877 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10878 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10879 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10880 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10881 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10882 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10883 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10884 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10885 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10886 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10887 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10888 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10889 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10890 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10891 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10892 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10893 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10894 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10895 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10896 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10897 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10898 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10899 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10900 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10901 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10902 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10903 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10904 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10905 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10906 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10907 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10908 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10909 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10910 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10911 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10912 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10913 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10914 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10915 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10916 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10917 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10918 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10919 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10920 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10921 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10922 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10923 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10924 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10925 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10926 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10927 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10928 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10929 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10930 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10931 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10932 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10933 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10934 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10935 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10936 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10937 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10938 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10939 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10940 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10941 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10942 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10943 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10944 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10945 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10946 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10947 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10948 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10949 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10950 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10951 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10952 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10953 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10954 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10955 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10956 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10957 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10958 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10959 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10960 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10961 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10962 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10963 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10964 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10965 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10966 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10967 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10968 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10969 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10970 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10971 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10972 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10973 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10974 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10975 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10976 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10977 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10978 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10979 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10980 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10981 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10982 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10983 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10984 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10985 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10986 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10987 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10988 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10989 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10990 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10991 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10992 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10993 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10994 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10995 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10996 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10997 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10998 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10999 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11000 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11001 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11002 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11003 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11004 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11005 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11006 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11007 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11008 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11009 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11010 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11011 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11012 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11013 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11014 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11015 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11016 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11017 tapered_buf_1/a_580_0# tapered_buf_1/a_160_n140# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11018 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11019 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11020 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11021 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11022 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11023 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11024 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11025 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11026 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11027 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11028 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11029 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11030 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11031 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11032 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11033 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11034 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11035 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11036 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11037 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11038 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11039 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11040 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11041 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11042 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11043 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11044 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11045 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11046 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11047 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11048 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11049 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11050 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11051 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11052 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11053 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11054 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11055 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11056 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11057 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11058 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11059 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11060 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11061 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11062 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11063 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11064 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11065 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11066 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11067 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11068 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11069 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11070 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11071 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11072 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11073 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11074 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11075 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11076 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11077 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11078 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11079 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11080 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11081 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11082 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11083 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11084 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11085 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11086 tapered_buf_1/a_160_n140# tapered_buf_1/in tapered_buf_1/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11087 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11088 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11089 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11090 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11091 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11092 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11093 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11094 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11095 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11096 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11097 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11098 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11099 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11100 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11101 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11102 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11103 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11104 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11105 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11106 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11107 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11108 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11109 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11110 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11111 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11112 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11113 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11114 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11115 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11116 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11117 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11118 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11119 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11120 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11121 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11122 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11123 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11124 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11125 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11126 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11127 tapered_buf_1/a_580_0# tapered_buf_1/a_160_n140# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11128 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11129 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11130 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11131 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11132 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11133 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11134 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11135 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11136 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11137 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11138 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11139 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11140 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11141 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11142 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11143 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11144 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11145 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11146 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11147 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11148 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11149 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11150 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11151 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11152 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11153 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11154 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11155 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11156 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11157 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11158 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11159 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11160 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11161 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11162 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11163 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11164 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11165 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11166 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11167 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11168 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11169 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11170 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11171 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11172 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11173 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11174 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11175 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11176 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11177 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11178 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11179 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11180 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11181 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11182 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11183 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11184 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11185 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11186 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11187 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11188 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11189 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11190 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11191 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11192 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11193 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11194 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11195 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11196 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11197 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11198 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11199 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11200 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11201 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11202 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11203 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11204 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11205 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11206 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11207 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11208 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11209 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11210 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11211 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11212 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11213 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11214 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11215 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11216 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11217 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11218 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11219 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11220 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11221 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11222 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11223 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11224 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11225 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11226 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11227 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11228 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11229 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11230 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11231 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11232 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11233 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11234 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11235 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11236 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11237 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11238 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11239 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11240 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11241 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11242 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11243 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11244 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11245 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11246 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11247 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11248 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11249 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11250 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11251 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11252 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11253 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11254 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11255 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11256 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11257 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11258 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11259 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11260 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11261 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11262 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11263 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11264 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11265 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11266 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11267 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11268 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11269 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11270 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11271 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11272 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11273 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11274 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11275 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11276 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11277 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11278 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11279 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11280 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11281 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11282 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11283 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11284 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11285 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11286 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11287 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11288 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11289 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11290 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11291 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11292 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11293 gnd tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11294 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11295 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11296 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11297 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11298 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11299 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11300 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11301 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11302 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11303 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11304 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11305 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11306 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11307 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11308 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11309 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11310 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11311 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11312 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11313 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11314 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11315 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11316 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11317 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11318 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11319 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11320 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11321 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11322 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11323 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11324 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11325 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11326 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11327 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11328 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11329 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11330 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11331 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11332 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11333 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11334 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11335 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11336 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11337 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11338 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11339 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11340 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11341 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11342 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11343 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11344 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11345 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11346 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11347 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11348 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11349 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11350 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11351 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11352 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11353 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11354 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11355 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11356 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11357 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11358 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11359 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11360 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11361 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11362 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11363 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11364 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11365 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11366 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11367 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11368 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11369 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11370 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11371 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11372 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11373 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11374 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11375 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11376 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11377 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11378 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11379 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11380 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11381 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11382 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11383 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11384 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11385 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11386 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11387 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11388 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11389 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11390 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11391 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11392 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11393 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11394 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11395 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11396 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11397 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11398 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11399 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11400 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11401 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11402 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11403 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11404 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11405 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11406 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11407 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11408 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11409 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11410 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11411 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11412 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11413 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11414 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11415 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11416 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11417 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11418 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11419 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11420 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11421 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11422 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11423 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11424 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11425 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11426 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11427 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11428 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11429 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11430 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11431 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11432 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11433 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11434 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11435 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11436 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11437 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11438 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11439 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11440 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11441 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11442 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11443 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11444 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11445 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11446 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11447 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11448 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11449 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11450 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11451 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11452 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11453 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11454 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11455 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11456 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11457 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11458 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11459 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11460 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11461 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11462 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11463 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11464 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11465 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11466 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11467 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11468 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11469 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11470 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11471 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11472 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11473 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11474 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11475 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11476 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11477 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11478 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11479 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11480 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11481 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11482 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11483 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11484 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11485 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11486 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11487 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11488 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11489 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11490 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11491 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11492 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11493 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11494 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11495 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11496 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11497 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11498 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11499 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11500 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11501 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11502 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11503 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11504 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11505 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11506 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11507 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11508 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11509 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11510 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11511 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11512 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11513 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11514 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11515 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11516 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11517 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11518 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11519 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11520 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11521 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11522 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11523 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11524 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11525 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11526 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11527 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11528 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11529 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11530 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11531 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11532 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11533 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11534 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11535 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11536 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11537 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11538 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11539 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11540 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11541 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11542 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11543 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11544 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11545 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11546 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11547 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11548 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11549 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11550 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11551 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11552 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11553 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11554 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11555 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11556 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11557 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11558 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11559 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11560 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11561 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11562 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11563 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11564 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11565 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11566 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11567 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11568 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11569 gnd tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11570 tapered_buf_1/a_580_0# tapered_buf_1/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11571 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11572 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11573 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11574 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11575 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11576 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11577 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11578 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11579 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11580 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11581 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11582 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11583 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11584 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11585 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11586 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11587 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11588 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11589 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11590 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11591 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11592 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11593 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11594 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11595 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11596 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11597 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11598 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11599 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11600 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11601 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11602 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11603 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11604 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11605 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11606 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11607 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11608 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11609 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11610 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11611 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11612 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11613 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11614 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11615 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11616 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11617 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11618 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11619 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11620 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11621 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11622 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11623 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11624 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11625 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11626 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11627 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11628 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11629 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11630 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11631 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11632 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11633 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11634 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11635 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11636 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11637 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11638 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11639 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11640 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11641 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11642 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11643 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11644 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11645 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11646 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11647 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11648 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11649 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11650 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11651 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11652 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11653 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11654 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11655 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11656 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11657 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11658 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11659 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11660 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11661 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11662 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11663 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11664 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11665 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11666 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11667 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11668 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11669 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11670 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11671 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11672 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11673 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11674 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11675 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11676 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11677 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11678 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11679 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11680 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11681 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11682 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11683 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11684 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11685 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11686 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11687 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11688 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11689 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11690 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11691 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11692 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11693 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11694 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11695 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11696 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11697 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11698 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11699 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11700 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11701 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11702 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11703 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11704 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11705 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11706 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11707 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11708 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11709 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11710 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11711 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11712 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11713 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11714 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11715 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11716 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11717 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11718 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11719 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11720 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11721 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11722 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11723 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11724 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11725 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11726 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11727 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11728 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11729 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11730 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11731 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11732 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11733 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11734 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11735 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11736 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11737 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11738 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11739 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11740 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11741 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11742 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11743 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11744 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11745 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11746 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11747 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11748 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11749 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11750 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11751 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11752 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11753 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11754 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11755 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11756 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11757 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11758 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11759 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11760 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11761 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11762 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11763 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11764 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11765 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11766 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11767 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11768 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11769 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11770 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11771 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11772 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11773 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11774 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11775 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11776 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11777 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11778 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11779 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11780 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11781 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11782 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11783 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11784 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11785 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11786 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11787 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11788 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11789 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11790 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11791 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11792 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11793 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11794 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11795 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11796 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11797 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11798 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11799 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11800 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11801 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11802 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11803 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11804 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11805 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11806 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11807 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11808 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11809 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11810 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11811 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11812 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11813 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11814 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11815 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11816 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11817 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11818 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11819 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11820 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11821 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11822 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11823 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11824 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11825 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11826 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11827 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11828 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11829 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11830 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11831 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11832 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11833 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11834 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11835 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11836 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11837 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11838 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11839 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11840 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11841 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11842 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11843 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11844 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11845 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11846 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11847 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11848 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11849 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11850 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11851 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11852 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11853 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11854 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11855 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11856 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11857 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11858 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11859 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11860 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11861 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11862 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11863 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11864 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11865 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11866 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11867 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11868 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11869 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11870 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11871 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11872 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11873 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11874 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11875 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11876 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11877 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11878 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11879 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11880 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11881 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11882 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11883 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11884 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11885 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11886 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11887 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11888 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11889 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11890 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11891 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11892 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11893 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11894 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11895 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11896 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11897 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11898 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11899 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11900 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11901 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11902 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11903 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11904 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11905 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11906 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11907 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11908 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11909 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11910 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11911 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11912 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11913 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11914 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11915 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11916 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11917 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11918 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11919 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11920 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11921 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11922 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11923 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11924 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11925 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11926 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11927 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11928 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11929 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11930 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11931 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11932 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11933 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11934 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11935 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11936 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11937 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11938 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11939 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11940 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11941 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11942 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11943 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11944 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11945 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11946 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11947 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11948 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11949 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11950 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11951 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11952 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11953 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11954 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11955 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11956 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11957 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11958 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11959 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11960 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11961 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11962 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11963 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11964 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11965 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11966 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11967 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11968 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11969 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11970 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11971 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11972 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11973 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11974 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11975 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11976 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11977 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11978 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11979 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11980 gnd tapered_buf_1/a_210_n610# tapered_buf_1/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11981 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11982 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11983 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11984 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11985 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11986 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11987 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11988 tapered_buf_1/out tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11989 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11990 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11991 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11992 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11993 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11994 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11995 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11996 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11997 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11998 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11999 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12000 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12001 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12002 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12003 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12004 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12005 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12006 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12007 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12008 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12009 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12010 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12011 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12012 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12013 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12014 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12015 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12016 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12017 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12018 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12019 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12020 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12021 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12022 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12023 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12024 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12025 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12026 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12027 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12028 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12029 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12030 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12031 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12032 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12033 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12034 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12035 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12036 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12037 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12038 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12039 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12040 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12041 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12042 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12043 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12044 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12045 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12046 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12047 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12048 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12049 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12050 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12051 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12052 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12053 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12054 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12055 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12056 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12057 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12058 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12059 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12060 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12061 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12062 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12063 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12064 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12065 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12066 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12067 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12068 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12069 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12070 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12071 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12072 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12073 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12074 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12075 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12076 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12077 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12078 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12079 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12080 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12081 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12082 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12083 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12084 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12085 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12086 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12087 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12088 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12089 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12090 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12091 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12092 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12093 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12094 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12095 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12096 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12097 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12098 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12099 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12100 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12101 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12102 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12103 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12104 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12105 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12106 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12107 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12108 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12109 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12110 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12111 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12112 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12113 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12114 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12115 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12116 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12117 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12118 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12119 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12120 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12121 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12122 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12123 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12124 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12125 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12126 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12127 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12128 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12129 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12130 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12131 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12132 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12133 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12134 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12135 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12136 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12137 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12138 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12139 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12140 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12141 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12142 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12143 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12144 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12145 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12146 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12147 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12148 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12149 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12150 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12151 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12152 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12153 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12154 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12155 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12156 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12157 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12158 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12159 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12160 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12161 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12162 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12163 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12164 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12165 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12166 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12167 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12168 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12169 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12170 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12171 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12172 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12173 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12174 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12175 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12176 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12177 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12178 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12179 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12180 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12181 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12182 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12183 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12184 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12185 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12186 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12187 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12188 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12189 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12190 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12191 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12192 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12193 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12194 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12195 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12196 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12197 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12198 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12199 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12200 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12201 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12202 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12203 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12204 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12205 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12206 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12207 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12208 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12209 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12210 tapered_buf_0/a_160_230# tapered_buf_0/in tapered_buf_0/a_n10_230# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12211 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12212 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12213 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12214 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12215 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12216 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12217 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12218 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12219 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12220 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12221 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12222 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12223 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12224 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12225 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12226 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12227 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12228 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12229 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12230 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12231 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12232 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12233 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12234 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12235 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12236 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12237 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12238 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12239 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12240 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12241 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12242 tapered_buf_0/a_580_0# tapered_buf_0/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12243 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12244 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12245 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12246 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12247 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12248 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12249 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12250 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12251 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12252 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12253 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12254 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12255 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12256 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12257 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12258 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12259 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12260 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12261 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12262 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12263 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12264 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12265 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12266 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12267 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12268 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12269 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12270 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12271 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12272 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12273 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12274 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12275 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12276 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12277 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12278 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12279 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12280 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12281 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12282 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12283 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12284 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12285 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12286 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12287 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12288 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12289 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12290 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12291 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12292 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12293 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12294 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12295 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12296 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12297 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12298 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12299 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12300 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12301 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12302 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12303 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12304 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12305 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12306 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12307 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12308 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12309 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12310 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12311 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12312 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12313 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12314 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12315 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12316 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12317 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12318 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12319 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12320 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12321 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12322 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12323 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12324 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12325 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12326 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12327 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12328 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12329 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12330 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12331 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12332 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12333 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12334 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12335 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12336 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12337 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12338 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12339 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12340 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12341 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12342 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12343 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12344 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12345 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12346 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12347 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12348 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12349 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12350 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12351 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12352 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12353 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12354 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12355 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12356 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12357 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12358 gnd tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12359 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12360 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12361 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12362 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12363 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12364 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12365 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12366 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12367 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12368 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12369 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12370 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12371 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12372 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12373 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12374 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12375 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12376 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12377 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12378 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12379 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12380 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12381 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12382 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12383 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12384 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12385 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12386 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12387 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12388 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12389 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12390 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12391 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12392 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12393 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12394 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12395 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12396 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12397 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12398 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12399 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12400 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12401 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12402 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12403 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12404 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12405 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12406 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12407 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12408 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12409 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12410 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12411 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12412 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12413 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12414 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12415 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12416 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12417 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12418 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12419 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12420 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12421 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12422 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12423 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12424 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12425 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12426 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12427 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12428 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12429 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12430 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12431 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12432 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12433 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12434 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12435 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12436 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12437 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12438 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12439 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12440 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12441 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12442 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12443 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12444 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12445 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12446 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12447 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12448 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12449 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12450 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12451 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12452 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12453 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12454 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12455 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12456 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12457 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12458 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12459 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12460 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12461 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12462 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12463 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12464 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12465 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12466 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12467 gnd tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12468 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12469 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12470 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12471 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12472 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12473 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12474 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12475 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12476 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12477 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12478 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12479 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12480 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12481 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12482 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12483 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12484 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12485 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12486 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12487 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12488 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12489 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12490 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12491 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12492 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12493 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12494 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12495 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12496 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12497 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12498 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12499 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12500 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12501 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12502 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12503 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12504 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12505 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12506 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12507 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12508 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12509 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12510 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12511 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12512 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12513 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12514 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12515 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12516 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12517 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12518 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12519 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12520 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12521 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12522 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12523 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12524 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12525 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12526 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12527 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12528 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12529 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12530 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12531 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12532 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12533 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12534 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12535 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12536 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12537 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12538 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12539 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12540 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12541 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12542 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12543 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12544 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12545 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12546 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12547 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12548 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12549 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12550 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12551 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12552 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12553 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12554 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12555 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12556 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12557 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12558 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12559 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12560 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12561 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12562 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12563 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12564 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12565 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12566 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12567 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12568 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12569 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12570 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12571 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12572 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12573 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12574 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12575 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12576 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12577 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12578 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12579 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12580 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12581 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12582 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12583 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12584 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12585 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12586 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12587 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12588 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12589 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12590 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12591 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12592 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12593 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12594 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12595 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12596 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12597 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12598 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12599 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12600 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12601 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12602 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12603 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12604 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12605 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12606 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12607 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12608 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12609 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12610 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12611 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12612 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12613 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12614 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12615 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12616 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12617 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12618 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12619 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12620 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12621 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12622 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12623 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12624 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12625 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12626 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12627 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12628 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12629 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12630 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12631 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12632 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12633 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12634 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12635 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12636 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12637 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12638 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12639 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12640 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12641 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12642 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12643 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12644 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12645 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12646 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12647 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12648 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12649 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12650 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12651 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12652 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12653 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12654 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12655 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12656 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12657 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12658 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12659 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12660 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12661 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12662 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12663 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12664 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12665 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12666 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12667 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12668 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12669 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12670 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12671 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12672 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12673 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12674 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12675 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12676 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12677 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12678 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12679 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12680 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12681 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12682 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12683 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12684 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12685 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12686 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12687 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12688 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12689 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12690 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12691 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12692 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12693 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12694 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12695 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12696 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12697 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12698 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12699 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12700 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12701 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12702 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12703 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12704 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12705 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12706 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12707 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12708 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12709 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12710 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12711 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12712 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12713 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12714 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12715 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12716 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12717 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12718 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12719 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12720 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12721 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12722 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12723 tapered_buf_0/a_580_0# tapered_buf_0/a_160_n140# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12724 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12725 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12726 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12727 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12728 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12729 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12730 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12731 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12732 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12733 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12734 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12735 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12736 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12737 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12738 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12739 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12740 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12741 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12742 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12743 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12744 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12745 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12746 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12747 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12748 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12749 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12750 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12751 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12752 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12753 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12754 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12755 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12756 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12757 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12758 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12759 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12760 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12761 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12762 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12763 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12764 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12765 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12766 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12767 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12768 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12769 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12770 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12771 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12772 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12773 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12774 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12775 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12776 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12777 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12778 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12779 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12780 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12781 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12782 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12783 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12784 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12785 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12786 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12787 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12788 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12789 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12790 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12791 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12792 tapered_buf_0/a_160_n140# tapered_buf_0/in tapered_buf_0/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12793 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12794 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12795 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12796 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12797 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12798 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12799 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12800 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12801 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12802 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12803 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12804 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12805 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12806 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12807 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12808 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12809 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12810 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12811 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12812 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12813 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12814 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12815 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12816 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12817 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12818 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12819 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12820 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12821 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12822 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12823 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12824 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12825 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12826 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12827 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12828 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12829 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12830 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12831 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12832 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12833 tapered_buf_0/a_580_0# tapered_buf_0/a_160_n140# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12834 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12835 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12836 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12837 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12838 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12839 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12840 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12841 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12842 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12843 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12844 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12845 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12846 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12847 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12848 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12849 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12850 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12851 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12852 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12853 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12854 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12855 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12856 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12857 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12858 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12859 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12860 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12861 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12862 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12863 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12864 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12865 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12866 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12867 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12868 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12869 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12870 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12871 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12872 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12873 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12874 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12875 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12876 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12877 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12878 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12879 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12880 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12881 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12882 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12883 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12884 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12885 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12886 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12887 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12888 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12889 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12890 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12891 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12892 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12893 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12894 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12895 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12896 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12897 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12898 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12899 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12900 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12901 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12902 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12903 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12904 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12905 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12906 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12907 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12908 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12909 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12910 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12911 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12912 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12913 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12914 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12915 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12916 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12917 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12918 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12919 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12920 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12921 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12922 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12923 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12924 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12925 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12926 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12927 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12928 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12929 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12930 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12931 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12932 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12933 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12934 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12935 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12936 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12937 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12938 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12939 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12940 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12941 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12942 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12943 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12944 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12945 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12946 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12947 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12948 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12949 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12950 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12951 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12952 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12953 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12954 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12955 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12956 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12957 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12958 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12959 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12960 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12961 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12962 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12963 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12964 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12965 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12966 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12967 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12968 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12969 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12970 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12971 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12972 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12973 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12974 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12975 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12976 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12977 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12978 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12979 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12980 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12981 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12982 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12983 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12984 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12985 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12986 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12987 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12988 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12989 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12990 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12991 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12992 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12993 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12994 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12995 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12996 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12997 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12998 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12999 gnd tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13000 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13001 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13002 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13003 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13004 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13005 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13006 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13007 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13008 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13009 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13010 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13011 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13012 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13013 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13014 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13015 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13016 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13017 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13018 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13019 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13020 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13021 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13022 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13023 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13024 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13025 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13026 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13027 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13028 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13029 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13030 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13031 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13032 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13033 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13034 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13035 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13036 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13037 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13038 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13039 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13040 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13041 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13042 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13043 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13044 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13045 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13046 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13047 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13048 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13049 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13050 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13051 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13052 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13053 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13054 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13055 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13056 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13057 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13058 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13059 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13060 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13061 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13062 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13063 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13064 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13065 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13066 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13067 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13068 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13069 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13070 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13071 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13072 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13073 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13074 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13075 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13076 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13077 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13078 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13079 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13080 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13081 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13082 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13083 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13084 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13085 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13086 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13087 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13088 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13089 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13090 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13091 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13092 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13093 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13094 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13095 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13096 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13097 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13098 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13099 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13100 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13101 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13102 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13103 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13104 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13105 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13106 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13107 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13108 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13109 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13110 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13111 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13112 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13113 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13114 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13115 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13116 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13117 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13118 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13119 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13120 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13121 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13122 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13123 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13124 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13125 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13126 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13127 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13128 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13129 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13130 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13131 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13132 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13133 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13134 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13135 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13136 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13137 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13138 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13139 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13140 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13141 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13142 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13143 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13144 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13145 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13146 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13147 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13148 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13149 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13150 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13151 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13152 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13153 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13154 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13155 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13156 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13157 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13158 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13159 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13160 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13161 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13162 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13163 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13164 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13165 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13166 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13167 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13168 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13169 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13170 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13171 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13172 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13173 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13174 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13175 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13176 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13177 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13178 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13179 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13180 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13181 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13182 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13183 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13184 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13185 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13186 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13187 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13188 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13189 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13190 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13191 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13192 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13193 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13194 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13195 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13196 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13197 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13198 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13199 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13200 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13201 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13202 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13203 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13204 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13205 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13206 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13207 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13208 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13209 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13210 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13211 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13212 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13213 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13214 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13215 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13216 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13217 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13218 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13219 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13220 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13221 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13222 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13223 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13224 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13225 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13226 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13227 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13228 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13229 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13230 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13231 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13232 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13233 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13234 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13235 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13236 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13237 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13238 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13239 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13240 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13241 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13242 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13243 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13244 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13245 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13246 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13247 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13248 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13249 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13250 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13251 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13252 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13253 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13254 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13255 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13256 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13257 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13258 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13259 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13260 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13261 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13262 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13263 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13264 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13265 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13266 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13267 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13268 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13269 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13270 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13271 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13272 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13273 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13274 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13275 gnd tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13276 tapered_buf_0/a_580_0# tapered_buf_0/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13277 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13278 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13279 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13280 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13281 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13282 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13283 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13284 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13285 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13286 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13287 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13288 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13289 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13290 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13291 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13292 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13293 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13294 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13295 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13296 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13297 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13298 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13299 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13300 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13301 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13302 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13303 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13304 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13305 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13306 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13307 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13308 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13309 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13310 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13311 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13312 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13313 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13314 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13315 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13316 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13317 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13318 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13319 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13320 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13321 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13322 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13323 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13324 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13325 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13326 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13327 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13328 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13329 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13330 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13331 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13332 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13333 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13334 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13335 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13336 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13337 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13338 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13339 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13340 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13341 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13342 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13343 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13344 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13345 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13346 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13347 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13348 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13349 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13350 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13351 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13352 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13353 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13354 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13355 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13356 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13357 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13358 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13359 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13360 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13361 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13362 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13363 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13364 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13365 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13366 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13367 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13368 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13369 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13370 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13371 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13372 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13373 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13374 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13375 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13376 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13377 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13378 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13379 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13380 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13381 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13382 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13383 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13384 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13385 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13386 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13387 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13388 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13389 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13390 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13391 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13392 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13393 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13394 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13395 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13396 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13397 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13398 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13399 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13400 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13401 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13402 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13403 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13404 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13405 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13406 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13407 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13408 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13409 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13410 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13411 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13412 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13413 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13414 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13415 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13416 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13417 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13418 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13419 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13420 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13421 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13422 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13423 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13424 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13425 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13426 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13427 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13428 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13429 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13430 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13431 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13432 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13433 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13434 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13435 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13436 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13437 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13438 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13439 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13440 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13441 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13442 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13443 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13444 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13445 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13446 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13447 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13448 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13449 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13450 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13451 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13452 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13453 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13454 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13455 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13456 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13457 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13458 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13459 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13460 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13461 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13462 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13463 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13464 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13465 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13466 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13467 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13468 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13469 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13470 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13471 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13472 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13473 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13474 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13475 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13476 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13477 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13478 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13479 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13480 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13481 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13482 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13483 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13484 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13485 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13486 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13487 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13488 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13489 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13490 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13491 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13492 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13493 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13494 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13495 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13496 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13497 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13498 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13499 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13500 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13501 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13502 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13503 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13504 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13505 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13506 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13507 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13508 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13509 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13510 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13511 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13512 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13513 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13514 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13515 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13516 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13517 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13518 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13519 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13520 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13521 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13522 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13523 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13524 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13525 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13526 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13527 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13528 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13529 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13530 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13531 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13532 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13533 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13534 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13535 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13536 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13537 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13538 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13539 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13540 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13541 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13542 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13543 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13544 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13545 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13546 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13547 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13548 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13549 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13550 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13551 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13552 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13553 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13554 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13555 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13556 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13557 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13558 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13559 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13560 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13561 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13562 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13563 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13564 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13565 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13566 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13567 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13568 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13569 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13570 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13571 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13572 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13573 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13574 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13575 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13576 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13577 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13578 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13579 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13580 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13581 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13582 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13583 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13584 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13585 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13586 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13587 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13588 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13589 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13590 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13591 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13592 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13593 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13594 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13595 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13596 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13597 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13598 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13599 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13600 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13601 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13602 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13603 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13604 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13605 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13606 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13607 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13608 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13609 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13610 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13611 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13612 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13613 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13614 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13615 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13616 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13617 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13618 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13619 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13620 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13621 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13622 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13623 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13624 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13625 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13626 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13627 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13628 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13629 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13630 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13631 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13632 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13633 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13634 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13635 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13636 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13637 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13638 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13639 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13640 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13641 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13642 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13643 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13644 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13645 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13646 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13647 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13648 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13649 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13650 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13651 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13652 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13653 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13654 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13655 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13656 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13657 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13658 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13659 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13660 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13661 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13662 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13663 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13664 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13665 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13666 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13667 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13668 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13669 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13670 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13671 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13672 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13673 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13674 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13675 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13676 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13677 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13678 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13679 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13680 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13681 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13682 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13683 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13684 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13685 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13686 gnd tapered_buf_0/a_210_n610# tapered_buf_0/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13687 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13688 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13689 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13690 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13691 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13692 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13693 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13694 tapered_buf_0/out tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13695 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
C0 tapered_buf_1/a_n10_n140# tapered_buf_1/a_160_n140# 0.05fF
C1 ro_complete_0/a4 ro_complete_0/cbank_1/v 0.05fF
C2 tapered_buf_4/a_n10_230# tapered_buf_4/a_n10_n140# 0.01fF
C3 tapered_buf_7/a_580_0# tapered_buf_7/a_160_230# 0.02fF
C4 ro_complete_0/a3 ro_complete_0/cbank_1/switch_4/vin 0.13fF
C5 ro_complete_0/cbank_0/switch_5/vin ro_complete_0/cbank_0/v 1.30fF
C6 ro_complete_0/cbank_0/switch_2/vin ro_complete_0/a2 0.09fF
C7 tapered_buf_5/a_160_n140# tapered_buf_5/a_210_n610# 0.22fF
C8 ro_complete_0/cbank_2/switch_1/vin ro_complete_0/cbank_2/switch_2/vin 0.20fF
C9 tapered_buf_3/a_580_0# tapered_buf_3/a_210_n610# 0.84fF
C10 tapered_buf_3/in tapered_buf_3/a_n10_n140# 0.04fF
C11 tapered_buf_6/a_160_n140# tapered_buf_6/a_580_0# 0.35fF
C12 ro_complete_0/a0 ro_complete_0/cbank_1/switch_1/vin 0.13fF
C13 tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# 4.78fF
C14 tapered_buf_1/a_n10_n140# tapered_buf_1/in 0.04fF
C15 tapered_buf_1/a_n10_230# tapered_buf_1/a_n10_n140# 0.01fF
C16 tapered_buf_1/in ro_complete_0/cbank_2/switch_0/vin 1.30fF
C17 tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# 1.27fF
C18 tapered_buf_2/in tapered_buf_2/a_n10_230# 0.02fF
C19 ro_complete_0/a3 ro_complete_0/a4 2.04fF
C20 ro_complete_0/a0 tapered_buf_1/in 0.05fF
C21 ro_complete_0/cbank_0/v tapered_buf_1/in 1.27fF
C22 tapered_buf_7/a_580_0# tapered_buf_7/a_210_n610# 0.84fF
C23 tapered_buf_7/in tapered_buf_7/a_n10_n140# 0.04fF
C24 tapered_buf_3/a_210_n610# ro_complete_0/a4 26.29fF
C25 tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# 0.35fF
C26 tapered_buf_5/a_1650_0# tapered_buf_5/a_210_n610# 2.89fF
C27 tapered_buf_5/a_n10_230# tapered_buf_5/a_160_230# 0.09fF
C28 tapered_buf_5/a_160_n140# tapered_buf_5/a_n10_n140# 0.05fF
C29 tapered_buf_7/a_210_n610# ro_complete_0/a0 26.29fF
C30 ro_complete_0/a2 ro_complete_0/cbank_2/switch_2/vin 0.09fF
C31 tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# 29.21fF
C32 tapered_buf_6/a_580_0# tapered_buf_6/a_1650_0# 1.27fF
C33 tapered_buf_6/in tapered_buf_6/a_n10_230# 0.02fF
C34 ro_complete_0/cbank_0/switch_1/vin ro_complete_0/cbank_0/switch_2/vin 0.20fF
C35 ro_complete_0/cbank_2/switch_1/vin ro_complete_0/cbank_2/switch_0/vin 0.20fF
C36 ro_complete_0/cbank_2/switch_4/vin tapered_buf_1/in 1.30fF
C37 ro_complete_0/a0 ro_complete_0/cbank_2/switch_1/vin 0.13fF
C38 tapered_buf_0/in tapered_buf_0/a_160_n140# 0.19fF
C39 ro_complete_0/cbank_0/switch_1/vin ro_complete_0/cbank_0/switch_0/vin 0.20fF
C40 tapered_buf_2/a_160_n140# tapered_buf_2/a_160_230# 0.17fF
C41 tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# 4.78fF
C42 ro_complete_0/a3 ro_complete_0/cbank_1/v 0.05fF
C43 ro_complete_0/cbank_2/switch_3/vin ro_complete_0/cbank_2/switch_4/vin 0.20fF
C44 tapered_buf_3/in tapered_buf_3/a_160_n140# 0.19fF
C45 ro_complete_0/a4 ro_complete_0/cbank_2/switch_5/vin 0.12fF
C46 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/a3 0.09fF
C47 tapered_buf_7/a_4670_0# tapered_buf_7/a_210_n610# 29.21fF
C48 tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# 1.27fF
C49 tapered_buf_5/a_210_n610# ro_complete_0/a2 26.29fF
C50 ro_complete_0/a1 ro_complete_0/cbank_1/v 0.05fF
C51 tapered_buf_6/a_160_n140# tapered_buf_6/a_160_230# 0.17fF
C52 tapered_buf_6/a_1650_0# tapered_buf_6/a_4670_0# 4.78fF
C53 tapered_buf_0/a_n10_n140# tapered_buf_0/a_160_n140# 0.05fF
C54 tapered_buf_1/a_160_n140# tapered_buf_1/in 0.19fF
C55 tapered_buf_4/a_580_0# tapered_buf_4/a_160_230# 0.02fF
C56 tapered_buf_7/in tapered_buf_7/a_160_n140# 0.19fF
C57 tapered_buf_2/a_160_n140# tapered_buf_2/a_210_n610# 0.22fF
C58 ro_complete_0/cbank_0/switch_5/vin ro_complete_0/a5 0.09fF
C59 tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# 0.35fF
C60 tapered_buf_1/a_210_n610# tapered_buf_1/a_160_n140# 0.22fF
C61 tapered_buf_1/a_n10_230# tapered_buf_1/in 0.02fF
C62 ro_complete_0/a0 ro_complete_0/cbank_1/switch_0/vin 0.09fF
C63 tapered_buf_5/a_n10_230# tapered_buf_5/a_n10_n140# 0.01fF
C64 ro_complete_0/cbank_2/switch_3/vin tapered_buf_1/in 1.30fF
C65 ro_complete_0/cbank_1/switch_5/vin ro_complete_0/a5 0.09fF
C66 tapered_buf_6/a_160_n140# tapered_buf_6/a_210_n610# 0.22fF
C67 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/cbank_0/switch_2/vin 0.20fF
C68 ro_complete_0/a5 tapered_buf_1/in 0.10fF
C69 tapered_buf_4/a_580_0# tapered_buf_4/a_210_n610# 0.84fF
C70 tapered_buf_4/in tapered_buf_4/a_n10_n140# 0.04fF
C71 tapered_buf_7/a_160_n140# tapered_buf_7/a_580_0# 0.35fF
C72 tapered_buf_0/a_160_230# tapered_buf_0/a_160_n140# 0.17fF
C73 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# 4.78fF
C74 tapered_buf_1/a_160_230# tapered_buf_1/a_580_0# 0.02fF
C75 tapered_buf_2/a_1650_0# tapered_buf_2/a_210_n610# 2.89fF
C76 tapered_buf_2/a_n10_230# tapered_buf_2/a_160_230# 0.09fF
C77 tapered_buf_2/a_160_n140# tapered_buf_2/a_n10_n140# 0.05fF
C78 tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# 1.27fF
C79 tapered_buf_3/in tapered_buf_3/a_n10_230# 0.02fF
C80 ro_complete_0/cbank_0/switch_1/vin ro_complete_0/a0 0.13fF
C81 ro_complete_0/cbank_2/switch_1/vin tapered_buf_1/in 1.30fF
C82 tapered_buf_0/in tapered_buf_0/a_n10_230# 0.02fF
C83 ro_complete_0/cbank_1/switch_1/vin ro_complete_0/cbank_1/switch_2/vin 0.20fF
C84 ro_complete_0/cbank_0/switch_1/vin ro_complete_0/cbank_0/v 1.30fF
C85 tapered_buf_0/a_580_0# tapered_buf_0/a_210_n610# 0.84fF
C86 ro_complete_0/cbank_0/switch_4/vin ro_complete_0/a4 0.09fF
C87 tapered_buf_6/a_1650_0# tapered_buf_6/a_210_n610# 2.89fF
C88 tapered_buf_6/a_n10_230# tapered_buf_6/a_160_230# 0.09fF
C89 tapered_buf_6/a_160_n140# tapered_buf_6/a_n10_n140# 0.05fF
C90 tapered_buf_4/a_4670_0# tapered_buf_4/a_210_n610# 29.21fF
C91 tapered_buf_7/a_580_0# tapered_buf_7/a_1650_0# 1.27fF
C92 tapered_buf_7/in tapered_buf_7/a_n10_230# 0.02fF
C93 tapered_buf_4/a_210_n610# ro_complete_0/a3 26.29fF
C94 ro_complete_0/cbank_0/switch_2/vin ro_complete_0/a1 0.14fF
C95 tapered_buf_3/a_160_n140# tapered_buf_3/a_160_230# 0.17fF
C96 tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# 4.78fF
C97 tapered_buf_0/a_n10_n140# tapered_buf_0/a_n10_230# 0.01fF
C98 ro_complete_0/a2 tapered_buf_1/in 0.05fF
C99 tapered_buf_4/in tapered_buf_4/a_160_n140# 0.19fF
C100 ro_complete_0/cbank_2/switch_3/vin ro_complete_0/a2 0.22fF
C101 tapered_buf_1/a_210_n610# tapered_buf_1/a_1650_0# 2.89fF
C102 ro_complete_0/cbank_1/switch_1/vin ro_complete_0/cbank_1/switch_0/vin 0.20fF
C103 ro_complete_0/a4 ro_complete_0/cbank_2/switch_4/vin 0.09fF
C104 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/cbank_0/switch_4/vin 0.20fF
C105 tapered_buf_7/a_160_n140# tapered_buf_7/a_160_230# 0.17fF
C106 tapered_buf_7/a_1650_0# tapered_buf_7/a_4670_0# 4.78fF
C107 tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# 29.21fF
C108 ro_complete_0/a0 ro_complete_0/cbank_1/v 0.05fF
C109 tapered_buf_2/a_n10_230# tapered_buf_2/a_n10_n140# 0.01fF
C110 tapered_buf_5/a_580_0# tapered_buf_5/a_160_230# 0.02fF
C111 ro_complete_0/a1 ro_complete_0/cbank_2/switch_2/vin 0.14fF
C112 ro_complete_0/cbank_0/v ro_complete_0/cbank_1/v 0.04fF
C113 tapered_buf_3/a_160_n140# tapered_buf_3/a_210_n610# 0.22fF
C114 tapered_buf_4/a_160_n140# tapered_buf_4/a_580_0# 0.35fF
C115 tapered_buf_0/a_n10_230# tapered_buf_0/a_160_230# 0.09fF
C116 ro_complete_0/cbank_0/switch_4/vin ro_complete_0/a3 0.13fF
C117 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/cbank_0/v 1.30fF
C118 ro_complete_0/cbank_0/switch_5/vin ro_complete_0/a4 0.12fF
C119 ro_complete_0/cbank_1/switch_4/vin ro_complete_0/cbank_1/switch_5/vin 0.19fF
C120 ro_complete_0/cbank_1/switch_2/vin ro_complete_0/a2 0.09fF
C121 tapered_buf_6/a_n10_230# tapered_buf_6/a_n10_n140# 0.01fF
C122 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/cbank_1/switch_2/vin 0.20fF
C123 tapered_buf_7/a_160_n140# tapered_buf_7/a_210_n610# 0.22fF
C124 tapered_buf_5/a_580_0# tapered_buf_5/a_210_n610# 0.84fF
C125 tapered_buf_5/in tapered_buf_5/a_n10_n140# 0.04fF
C126 ro_complete_0/cbank_1/switch_5/vin ro_complete_0/a4 0.12fF
C127 tapered_buf_3/a_1650_0# tapered_buf_3/a_210_n610# 2.89fF
C128 tapered_buf_3/a_n10_230# tapered_buf_3/a_160_230# 0.09fF
C129 tapered_buf_3/a_160_n140# tapered_buf_3/a_n10_n140# 0.05fF
C130 ro_complete_0/a4 tapered_buf_1/in 0.05fF
C131 tapered_buf_4/a_580_0# tapered_buf_4/a_1650_0# 1.27fF
C132 tapered_buf_4/in tapered_buf_4/a_n10_230# 0.02fF
C133 ro_complete_0/a0 ro_complete_0/a1 3.46fF
C134 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/a2 0.14fF
C135 ro_complete_0/a3 ro_complete_0/cbank_2/switch_4/vin 0.13fF
C136 ro_complete_0/a4 ro_complete_0/a5 2.39fF
C137 tapered_buf_7/a_1650_0# tapered_buf_7/a_210_n610# 2.89fF
C138 tapered_buf_7/a_n10_230# tapered_buf_7/a_160_230# 0.09fF
C139 tapered_buf_7/a_160_n140# tapered_buf_7/a_n10_n140# 0.05fF
C140 ro_complete_0/cbank_1/switch_1/vin ro_complete_0/cbank_1/v 1.30fF
C141 tapered_buf_5/a_4670_0# tapered_buf_5/a_210_n610# 29.21fF
C142 ro_complete_0/cbank_1/switch_5/vin ro_complete_0/cbank_1/v 1.45fF
C143 tapered_buf_1/out tapered_buf_1/a_210_n610# 26.29fF
C144 ro_complete_0/cbank_1/v tapered_buf_1/in 1.36fF
C145 tapered_buf_4/a_160_n140# tapered_buf_4/a_160_230# 0.17fF
C146 tapered_buf_4/a_1650_0# tapered_buf_4/a_4670_0# 4.78fF
C147 tapered_buf_2/a_210_n610# ro_complete_0/a5 26.29fF
C148 ro_complete_0/cbank_0/switch_2/vin ro_complete_0/cbank_0/v 1.30fF
C149 ro_complete_0/a0 ro_complete_0/cbank_0/switch_0/vin 0.09fF
C150 tapered_buf_2/a_580_0# tapered_buf_2/a_160_230# 0.02fF
C151 tapered_buf_5/in tapered_buf_5/a_160_n140# 0.19fF
C152 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_0/vin 1.30fF
C153 tapered_buf_6/a_210_n610# ro_complete_0/a1 26.29fF
C154 tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# 0.35fF
C155 ro_complete_0/cbank_1/v ro_complete_0/a5 0.08fF
C156 ro_complete_0/cbank_2/switch_4/vin ro_complete_0/cbank_2/switch_5/vin 0.19fF
C157 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/cbank_1/switch_4/vin 0.20fF
C158 ro_complete_0/a3 tapered_buf_1/in 0.05fF
C159 tapered_buf_3/a_n10_230# tapered_buf_3/a_n10_n140# 0.01fF
C160 tapered_buf_6/a_580_0# tapered_buf_6/a_160_230# 0.02fF
C161 tapered_buf_4/a_160_n140# tapered_buf_4/a_210_n610# 0.22fF
C162 tapered_buf_1/a_160_230# tapered_buf_1/a_160_n140# 0.17fF
C163 ro_complete_0/a3 ro_complete_0/cbank_2/switch_3/vin 0.21fF
C164 tapered_buf_2/a_580_0# tapered_buf_2/a_210_n610# 0.84fF
C165 tapered_buf_2/in tapered_buf_2/a_n10_n140# 0.04fF
C166 tapered_buf_5/a_160_n140# tapered_buf_5/a_580_0# 0.35fF
C167 ro_complete_0/cbank_1/switch_2/vin ro_complete_0/cbank_1/v 1.30fF
C168 tapered_buf_0/a_n10_n140# tapered_buf_0/in 0.04fF
C169 ro_complete_0/a1 tapered_buf_1/in 0.05fF
C170 tapered_buf_7/a_n10_230# tapered_buf_7/a_n10_n140# 0.01fF
C171 tapered_buf_0/a_160_n140# tapered_buf_0/a_210_n610# 0.22fF
C172 tapered_buf_1/a_210_n610# tapered_buf_1/a_580_0# 0.84fF
C173 tapered_buf_1/a_n10_230# tapered_buf_1/a_160_230# 0.09fF
C174 ro_complete_0/a2 ro_complete_0/cbank_1/v 0.05fF
C175 tapered_buf_6/a_580_0# tapered_buf_6/a_210_n610# 0.84fF
C176 tapered_buf_6/in tapered_buf_6/a_n10_n140# 0.04fF
C177 ro_complete_0/cbank_2/switch_5/vin tapered_buf_1/in 1.43fF
C178 tapered_buf_4/a_1650_0# tapered_buf_4/a_210_n610# 2.89fF
C179 tapered_buf_4/a_n10_230# tapered_buf_4/a_160_230# 0.09fF
C180 tapered_buf_4/a_160_n140# tapered_buf_4/a_n10_n140# 0.05fF
C181 tapered_buf_0/a_160_230# tapered_buf_0/a_580_0# 0.02fF
C182 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/a2 0.14fF
C183 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/cbank_1/v 1.30fF
C184 ro_complete_0/cbank_0/switch_4/vin ro_complete_0/cbank_0/v 1.30fF
C185 tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# 29.21fF
C186 tapered_buf_5/a_580_0# tapered_buf_5/a_1650_0# 1.27fF
C187 tapered_buf_5/in tapered_buf_5/a_n10_230# 0.02fF
C188 ro_complete_0/a1 ro_complete_0/cbank_2/switch_1/vin 0.14fF
C189 ro_complete_0/a0 ro_complete_0/cbank_2/switch_0/vin 0.09fF
C190 ro_complete_0/cbank_1/switch_4/vin ro_complete_0/a4 0.09fF
C191 tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# 1.27fF
C192 ro_complete_0/a5 ro_complete_0/cbank_2/switch_5/vin 0.09fF
C193 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_0/vin 1.30fF
C194 tapered_buf_2/in tapered_buf_2/a_160_n140# 0.19fF
C195 ro_complete_0/a3 ro_complete_0/a2 3.17fF
C196 tapered_buf_0/a_1650_0# tapered_buf_0/a_210_n610# 2.89fF
C197 ro_complete_0/cbank_1/switch_2/vin ro_complete_0/a1 0.14fF
C198 tapered_buf_6/a_4670_0# tapered_buf_6/a_210_n610# 29.21fF
C199 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/a3 0.09fF
C200 tapered_buf_5/a_160_n140# tapered_buf_5/a_160_230# 0.17fF
C201 tapered_buf_5/a_1650_0# tapered_buf_5/a_4670_0# 4.78fF
C202 ro_complete_0/a1 ro_complete_0/a2 3.18fF
C203 ro_complete_0/cbank_1/switch_4/vin ro_complete_0/cbank_1/v 1.30fF
C204 tapered_buf_3/a_580_0# tapered_buf_3/a_160_230# 0.02fF
C205 tapered_buf_6/in tapered_buf_6/a_160_n140# 0.19fF
C206 ro_complete_0/cbank_2/switch_2/vin tapered_buf_1/in 1.30fF
C207 ro_complete_0/cbank_0/switch_4/vin ro_complete_0/cbank_0/switch_5/vin 0.19fF
C208 tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# 0.35fF
C209 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# 29.21fF
C210 ro_complete_0/cbank_2/switch_3/vin ro_complete_0/cbank_2/switch_2/vin 0.20fF
C211 tapered_buf_0/a_n10_n140# tapered_buf_0/w_70_n1420# 0.06fF
C212 tapered_buf_0/a_210_n610# tapered_buf_0/w_70_n1420# 614.83fF
C213 tapered_buf_0/a_160_230# tapered_buf_0/w_70_n1420# 0.15fF
C214 tapered_buf_0/a_n10_230# tapered_buf_0/w_70_n1420# 0.13fF
C215 tapered_buf_0/a_4670_0# tapered_buf_0/w_70_n1420# 250.63fF
C216 tapered_buf_0/a_1650_0# tapered_buf_0/w_70_n1420# 63.04fF
C217 tapered_buf_0/a_580_0# tapered_buf_0/w_70_n1420# 16.64fF
C218 tapered_buf_0/a_160_n140# tapered_buf_0/w_70_n1420# 4.00fF
C219 tapered_buf_0/in tapered_buf_0/w_70_n1420# 1.13fF
C220 tapered_buf_1/out tapered_buf_0/w_70_n1420# 385.11fF
C221 tapered_buf_1/a_n10_n140# tapered_buf_0/w_70_n1420# 0.06fF
C222 tapered_buf_1/a_210_n610# tapered_buf_0/w_70_n1420# 588.54fF
C223 tapered_buf_1/a_160_230# tapered_buf_0/w_70_n1420# 0.15fF
C224 tapered_buf_1/a_n10_230# tapered_buf_0/w_70_n1420# 0.13fF
C225 tapered_buf_1/a_4670_0# tapered_buf_0/w_70_n1420# 250.63fF
C226 tapered_buf_1/a_1650_0# tapered_buf_0/w_70_n1420# 63.04fF
C227 tapered_buf_1/a_580_0# tapered_buf_0/w_70_n1420# 16.64fF
C228 tapered_buf_1/a_160_n140# tapered_buf_0/w_70_n1420# 4.00fF
C229 ro_complete_0/cbank_2/switch_0/vin tapered_buf_0/w_70_n1420# 1.30fF
C230 tapered_buf_1/in tapered_buf_0/w_70_n1420# 23.92fF
C231 ro_complete_0/cbank_2/switch_5/vin tapered_buf_0/w_70_n1420# 1.06fF
C232 ro_complete_0/a5 tapered_buf_0/w_70_n1420# 400.71fF
C233 ro_complete_0/cbank_2/switch_4/vin tapered_buf_0/w_70_n1420# 1.16fF
C234 ro_complete_0/a4 tapered_buf_0/w_70_n1420# 401.22fF
C235 ro_complete_0/cbank_2/switch_2/vin tapered_buf_0/w_70_n1420# 0.95fF
C236 ro_complete_0/a2 tapered_buf_0/w_70_n1420# 408.04fF
C237 ro_complete_0/cbank_2/switch_3/vin tapered_buf_0/w_70_n1420# 1.30fF
C238 ro_complete_0/a3 tapered_buf_0/w_70_n1420# 404.01fF
C239 ro_complete_0/cbank_2/switch_1/vin tapered_buf_0/w_70_n1420# 1.53fF
C240 ro_complete_0/a1 tapered_buf_0/w_70_n1420# 411.87fF
C241 ro_complete_0/a0 tapered_buf_0/w_70_n1420# 415.94fF
C242 ro_complete_0/cbank_1/switch_0/vin tapered_buf_0/w_70_n1420# 1.30fF
C243 ro_complete_0/cbank_1/v tapered_buf_0/w_70_n1420# 17.28fF
C244 ro_complete_0/cbank_1/switch_5/vin tapered_buf_0/w_70_n1420# 1.06fF
C245 ro_complete_0/cbank_1/switch_4/vin tapered_buf_0/w_70_n1420# 1.16fF
C246 ro_complete_0/cbank_1/switch_2/vin tapered_buf_0/w_70_n1420# 0.95fF
C247 ro_complete_0/cbank_1/switch_3/vin tapered_buf_0/w_70_n1420# 1.30fF
C248 ro_complete_0/cbank_1/switch_1/vin tapered_buf_0/w_70_n1420# 1.53fF
C249 ro_complete_0/cbank_0/switch_0/vin tapered_buf_0/w_70_n1420# 1.30fF
C250 ro_complete_0/cbank_0/v tapered_buf_0/w_70_n1420# 15.10fF
C251 ro_complete_0/cbank_0/switch_5/vin tapered_buf_0/w_70_n1420# 1.06fF
C252 ro_complete_0/cbank_0/switch_4/vin tapered_buf_0/w_70_n1420# 1.16fF
C253 ro_complete_0/cbank_0/switch_2/vin tapered_buf_0/w_70_n1420# 0.95fF
C254 ro_complete_0/cbank_0/switch_3/vin tapered_buf_0/w_70_n1420# 1.30fF
C255 ro_complete_0/cbank_0/switch_1/vin tapered_buf_0/w_70_n1420# 1.53fF
C256 tapered_buf_7/a_n10_n140# tapered_buf_0/w_70_n1420# 0.06fF
C257 tapered_buf_7/a_210_n610# tapered_buf_0/w_70_n1420# 588.54fF
C258 tapered_buf_7/a_160_230# tapered_buf_0/w_70_n1420# 0.15fF
C259 tapered_buf_7/a_n10_230# tapered_buf_0/w_70_n1420# 0.13fF
C260 tapered_buf_7/a_4670_0# tapered_buf_0/w_70_n1420# 250.63fF
C261 tapered_buf_7/a_1650_0# tapered_buf_0/w_70_n1420# 63.04fF
C262 tapered_buf_7/a_580_0# tapered_buf_0/w_70_n1420# 16.64fF
C263 tapered_buf_7/a_160_n140# tapered_buf_0/w_70_n1420# 4.00fF
C264 tapered_buf_7/in tapered_buf_0/w_70_n1420# 1.13fF
C265 tapered_buf_6/a_n10_n140# tapered_buf_0/w_70_n1420# 0.06fF
C266 tapered_buf_6/a_210_n610# tapered_buf_0/w_70_n1420# 588.54fF
C267 tapered_buf_6/a_160_230# tapered_buf_0/w_70_n1420# 0.15fF
C268 tapered_buf_6/a_n10_230# tapered_buf_0/w_70_n1420# 0.13fF
C269 tapered_buf_6/a_4670_0# tapered_buf_0/w_70_n1420# 250.63fF
C270 tapered_buf_6/a_1650_0# tapered_buf_0/w_70_n1420# 63.04fF
C271 tapered_buf_6/a_580_0# tapered_buf_0/w_70_n1420# 16.64fF
C272 tapered_buf_6/a_160_n140# tapered_buf_0/w_70_n1420# 4.00fF
C273 tapered_buf_6/in tapered_buf_0/w_70_n1420# 1.13fF
C274 tapered_buf_5/a_n10_n140# tapered_buf_0/w_70_n1420# 0.06fF
C275 tapered_buf_5/a_210_n610# tapered_buf_0/w_70_n1420# 588.54fF
C276 tapered_buf_5/a_160_230# tapered_buf_0/w_70_n1420# 0.15fF
C277 tapered_buf_5/a_n10_230# tapered_buf_0/w_70_n1420# 0.13fF
C278 tapered_buf_5/a_4670_0# tapered_buf_0/w_70_n1420# 250.63fF
C279 tapered_buf_5/a_1650_0# tapered_buf_0/w_70_n1420# 63.04fF
C280 tapered_buf_5/a_580_0# tapered_buf_0/w_70_n1420# 16.64fF
C281 tapered_buf_5/a_160_n140# tapered_buf_0/w_70_n1420# 4.00fF
C282 tapered_buf_5/in tapered_buf_0/w_70_n1420# 1.13fF
C283 tapered_buf_4/a_n10_n140# tapered_buf_0/w_70_n1420# 0.06fF
C284 tapered_buf_4/a_210_n610# tapered_buf_0/w_70_n1420# 588.54fF
C285 tapered_buf_4/a_160_230# tapered_buf_0/w_70_n1420# 0.15fF
C286 tapered_buf_4/a_n10_230# tapered_buf_0/w_70_n1420# 0.13fF
C287 tapered_buf_4/a_4670_0# tapered_buf_0/w_70_n1420# 250.63fF
C288 tapered_buf_4/a_1650_0# tapered_buf_0/w_70_n1420# 63.04fF
C289 tapered_buf_4/a_580_0# tapered_buf_0/w_70_n1420# 16.64fF
C290 tapered_buf_4/a_160_n140# tapered_buf_0/w_70_n1420# 4.00fF
C291 tapered_buf_4/in tapered_buf_0/w_70_n1420# 1.13fF
C292 tapered_buf_3/a_n10_n140# tapered_buf_0/w_70_n1420# 0.06fF
C293 tapered_buf_3/a_210_n610# tapered_buf_0/w_70_n1420# 588.54fF
C294 tapered_buf_3/a_160_230# tapered_buf_0/w_70_n1420# 0.15fF
C295 tapered_buf_3/a_n10_230# tapered_buf_0/w_70_n1420# 0.13fF
C296 tapered_buf_3/a_4670_0# tapered_buf_0/w_70_n1420# 250.63fF
C297 tapered_buf_3/a_1650_0# tapered_buf_0/w_70_n1420# 63.04fF
C298 tapered_buf_3/a_580_0# tapered_buf_0/w_70_n1420# 16.64fF
C299 tapered_buf_3/a_160_n140# tapered_buf_0/w_70_n1420# 4.00fF
C300 tapered_buf_3/in tapered_buf_0/w_70_n1420# 1.13fF
C301 tapered_buf_2/a_n10_n140# tapered_buf_0/w_70_n1420# 0.06fF
C302 tapered_buf_2/a_210_n610# tapered_buf_0/w_70_n1420# 588.54fF
C303 tapered_buf_2/a_160_230# tapered_buf_0/w_70_n1420# 0.15fF
C304 tapered_buf_2/a_n10_230# tapered_buf_0/w_70_n1420# 0.13fF
C305 tapered_buf_2/a_4670_0# tapered_buf_0/w_70_n1420# 250.63fF
C306 tapered_buf_2/a_1650_0# tapered_buf_0/w_70_n1420# 63.04fF
C307 tapered_buf_2/a_580_0# tapered_buf_0/w_70_n1420# 16.64fF
C308 tapered_buf_2/a_160_n140# tapered_buf_0/w_70_n1420# 4.00fF
C309 tapered_buf_2/in tapered_buf_0/w_70_n1420# 1.13fF

.ic v(out) 0
.tran 0.01ns 100ns

.control
run
  set hcopypscolor = 1
  set color0=white
  set color1=black

  hardcopy plots/ro_post.eps v(out)
.endc
.end