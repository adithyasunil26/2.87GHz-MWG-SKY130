magic
tech sky130A
timestamp 1713075058
<< psubdiff >>
rect 132 -121 262 -106
rect 132 -221 147 -121
rect 247 -221 262 -121
rect 132 -236 262 -221
rect 4121 -337 4251 -322
rect 4121 -437 4136 -337
rect 4236 -437 4251 -337
rect 4121 -452 4251 -437
rect 132 -611 262 -596
rect 132 -711 147 -611
rect 247 -711 262 -611
rect 132 -726 262 -711
rect 4121 -923 4251 -908
rect 4121 -1023 4136 -923
rect 4236 -1023 4251 -923
rect 4121 -1038 4251 -1023
rect 132 -1101 262 -1086
rect 132 -1201 147 -1101
rect 247 -1201 262 -1101
rect 132 -1216 262 -1201
rect 132 -1458 262 -1443
rect 132 -1558 147 -1458
rect 247 -1558 262 -1458
rect 132 -1573 262 -1558
rect 132 -1948 262 -1933
rect 132 -2048 147 -1948
rect 247 -2048 262 -1948
rect 132 -2063 262 -2048
rect 4121 -2329 4251 -2314
rect 132 -2438 262 -2423
rect 132 -2538 147 -2438
rect 247 -2538 262 -2438
rect 4121 -2429 4136 -2329
rect 4236 -2429 4251 -2329
rect 4121 -2444 4251 -2429
rect 132 -2553 262 -2538
rect 132 -2803 262 -2788
rect 132 -2903 147 -2803
rect 247 -2903 262 -2803
rect 132 -2918 262 -2903
rect 4121 -3149 4251 -3134
rect 4121 -3249 4136 -3149
rect 4236 -3249 4251 -3149
rect 4121 -3264 4251 -3249
rect 132 -3293 262 -3278
rect 132 -3393 147 -3293
rect 247 -3393 262 -3293
rect 132 -3408 262 -3393
rect 132 -3783 262 -3768
rect 132 -3883 147 -3783
rect 247 -3883 262 -3783
rect 132 -3898 262 -3883
rect 4146 -3949 4251 -3948
rect 4121 -3963 4251 -3949
rect 4121 -4063 4136 -3963
rect 4236 -4063 4251 -3963
rect 4121 -4078 4251 -4063
rect 132 -4148 262 -4133
rect 132 -4248 147 -4148
rect 247 -4248 262 -4148
rect 132 -4263 262 -4248
rect 4121 -4437 4251 -4422
rect 4121 -4537 4136 -4437
rect 4236 -4537 4251 -4437
rect 4121 -4552 4251 -4537
rect 132 -4638 262 -4623
rect 132 -4738 147 -4638
rect 247 -4738 262 -4638
rect 132 -4753 262 -4738
rect 4121 -5023 4251 -5008
rect 132 -5128 262 -5113
rect 132 -5228 147 -5128
rect 247 -5228 262 -5128
rect 4121 -5123 4136 -5023
rect 4236 -5123 4251 -5023
rect 4121 -5138 4251 -5123
rect 132 -5243 262 -5228
rect 560 -5562 690 -5547
rect 560 -5662 575 -5562
rect 675 -5662 690 -5562
rect 560 -5677 690 -5662
rect 1076 -5569 1206 -5554
rect 1076 -5669 1091 -5569
rect 1191 -5669 1206 -5569
rect 1076 -5684 1206 -5669
rect 1730 -5565 1860 -5550
rect 1730 -5665 1745 -5565
rect 1845 -5665 1860 -5565
rect 1730 -5680 1860 -5665
rect 2382 -5565 2512 -5550
rect 2382 -5665 2397 -5565
rect 2497 -5665 2512 -5565
rect 2382 -5680 2512 -5665
rect 3034 -5565 3164 -5550
rect 3034 -5665 3049 -5565
rect 3149 -5665 3164 -5565
rect 3034 -5680 3164 -5665
rect 3780 -5565 3910 -5550
rect 3780 -5665 3795 -5565
rect 3895 -5665 3910 -5565
rect 3780 -5680 3910 -5665
<< psubdiffcont >>
rect 147 -221 247 -121
rect 4136 -437 4236 -337
rect 147 -711 247 -611
rect 4136 -1023 4236 -923
rect 147 -1201 247 -1101
rect 147 -1558 247 -1458
rect 147 -2048 247 -1948
rect 147 -2538 247 -2438
rect 4136 -2429 4236 -2329
rect 147 -2903 247 -2803
rect 4136 -3249 4236 -3149
rect 147 -3393 247 -3293
rect 147 -3883 247 -3783
rect 4136 -4063 4236 -3963
rect 147 -4248 247 -4148
rect 4136 -4537 4236 -4437
rect 147 -4738 247 -4638
rect 147 -5228 247 -5128
rect 4136 -5123 4236 -5023
rect 575 -5662 675 -5562
rect 1091 -5669 1191 -5569
rect 1745 -5665 1845 -5565
rect 2397 -5665 2497 -5565
rect 3049 -5665 3149 -5565
rect 3795 -5665 3895 -5565
<< locali >>
rect 3720 750 3810 760
rect 665 740 735 750
rect 665 730 675 740
rect 505 700 675 730
rect 665 690 675 700
rect 725 690 735 740
rect 2210 735 2280 745
rect 2210 725 2220 735
rect 2040 695 2220 725
rect 665 680 735 690
rect 2210 685 2220 695
rect 2270 685 2280 735
rect 3720 730 3730 750
rect 3570 700 3730 730
rect 2210 675 2280 685
rect 3720 680 3730 700
rect 3800 680 3810 750
rect 3720 670 3810 680
rect 3598 420 3628 426
rect 3598 415 3632 420
rect 3598 338 3606 415
rect 3623 338 3632 415
rect 3598 336 3632 338
rect 3598 330 3628 336
rect 115 81 300 245
rect 4111 132 4261 147
rect 115 -121 275 81
rect 4108 -42 4266 132
rect 115 -221 147 -121
rect 247 -221 275 -121
rect 115 -611 275 -221
rect 115 -711 147 -611
rect 247 -711 275 -611
rect 115 -1101 275 -711
rect 4111 -337 4261 -42
rect 4111 -437 4136 -337
rect 4236 -437 4261 -337
rect 958 -840 1143 -805
rect 1462 -840 1632 -805
rect 1936 -840 2121 -805
rect 2426 -840 2606 -805
rect 2917 -840 3097 -805
rect 3428 -840 3693 -805
rect 115 -1201 147 -1101
rect 247 -1201 275 -1101
rect 115 -1458 275 -1201
rect 115 -1558 147 -1458
rect 247 -1558 275 -1458
rect 115 -1634 275 -1558
rect 425 -1634 981 -1633
rect 115 -1763 981 -1634
rect 115 -1764 565 -1763
rect 115 -1948 275 -1764
rect 115 -2048 147 -1948
rect 247 -2048 275 -1948
rect 115 -2438 275 -2048
rect 115 -2538 147 -2438
rect 247 -2538 275 -2438
rect 115 -2803 275 -2538
rect 1108 -2575 1143 -840
rect 1597 -2575 1632 -840
rect 2086 -2575 2121 -840
rect 2571 -2575 2606 -840
rect 3062 -2575 3097 -840
rect 3658 -2575 3693 -840
rect 4111 -923 4261 -437
rect 4111 -1023 4136 -923
rect 4236 -1023 4261 -923
rect 4111 -1468 4261 -1023
rect 4108 -1826 4264 -1468
rect 958 -2610 1143 -2575
rect 1462 -2610 1632 -2575
rect 1936 -2610 2121 -2575
rect 2426 -2610 2606 -2575
rect 2917 -2610 3097 -2575
rect 3428 -2610 3693 -2575
rect 115 -2903 147 -2803
rect 247 -2903 275 -2803
rect 115 -3293 275 -2903
rect 115 -3393 147 -3293
rect 247 -3393 275 -3293
rect 115 -3404 275 -3393
rect 382 -3404 967 -3401
rect 115 -3533 967 -3404
rect 115 -3534 563 -3533
rect 115 -3783 275 -3534
rect 115 -3883 147 -3783
rect 247 -3883 275 -3783
rect 115 -4148 275 -3883
rect 115 -4248 147 -4148
rect 247 -4248 275 -4148
rect 115 -4638 275 -4248
rect 1108 -4360 1143 -2610
rect 1597 -4360 1632 -2610
rect 2086 -4360 2121 -2610
rect 2571 -4360 2606 -2610
rect 3062 -4360 3097 -2610
rect 3658 -3649 3693 -2610
rect 4111 -2329 4261 -1826
rect 4111 -2429 4136 -2329
rect 4236 -2429 4261 -2329
rect 4111 -3149 4261 -2429
rect 4111 -3238 4136 -3149
rect 4108 -3249 4136 -3238
rect 4236 -3249 4261 -3149
rect 4108 -3598 4261 -3249
rect 3657 -3857 3694 -3649
rect 3658 -4360 3693 -3857
rect 958 -4395 1143 -4360
rect 1462 -4395 1632 -4360
rect 1936 -4395 2121 -4360
rect 2426 -4395 2606 -4360
rect 2917 -4395 3097 -4360
rect 3428 -4395 3693 -4360
rect 4111 -3963 4261 -3598
rect 4111 -4063 4136 -3963
rect 4236 -4063 4261 -3963
rect 115 -4738 147 -4638
rect 247 -4738 275 -4638
rect 115 -5128 275 -4738
rect 115 -5228 147 -5128
rect 247 -5191 275 -5128
rect 4111 -4437 4261 -4063
rect 4111 -4537 4136 -4437
rect 4236 -4537 4261 -4437
rect 4111 -5023 4261 -4537
rect 4111 -5123 4136 -5023
rect 4236 -5123 4261 -5023
rect 4111 -5136 4261 -5123
rect 406 -5191 991 -5190
rect 247 -5228 991 -5191
rect 115 -5318 991 -5228
rect 113 -5321 991 -5318
rect 113 -5528 276 -5321
rect 406 -5322 991 -5321
rect 4105 -5423 4261 -5136
rect 4105 -5426 4263 -5423
rect 4110 -5525 4263 -5426
rect 113 -5530 529 -5528
rect 663 -5530 4263 -5525
rect 113 -5562 4263 -5530
rect 113 -5662 575 -5562
rect 675 -5565 4263 -5562
rect 675 -5569 1745 -5565
rect 675 -5662 1091 -5569
rect 113 -5669 1091 -5662
rect 1191 -5665 1745 -5569
rect 1845 -5665 2397 -5565
rect 2497 -5665 3049 -5565
rect 3149 -5665 3795 -5565
rect 3895 -5665 4263 -5565
rect 1191 -5669 4263 -5665
rect 113 -5688 4263 -5669
rect 113 -5690 529 -5688
rect 663 -5693 4263 -5688
<< viali >>
rect 675 690 725 740
rect 2220 685 2270 735
rect 3730 680 3800 750
rect 3606 338 3623 415
<< metal1 >>
rect 3720 750 3810 760
rect 665 740 735 750
rect 665 690 675 740
rect 725 690 735 740
rect 665 680 735 690
rect 2210 735 2280 745
rect 2210 685 2220 735
rect 2270 685 2280 735
rect 2210 675 2280 685
rect 3720 680 3730 750
rect 3800 680 3810 750
rect 3720 670 3810 680
rect 3598 415 3628 426
rect 675 371 725 372
rect 3598 338 3606 415
rect 3623 338 3628 415
rect 3598 330 3628 338
<< via1 >>
rect 675 690 725 740
rect 2220 685 2270 735
rect 3730 680 3800 750
<< metal2 >>
rect 3710 750 4120 775
rect 665 740 735 750
rect 665 690 675 740
rect 725 690 735 740
rect 665 680 735 690
rect 2210 735 2280 745
rect 2210 685 2220 735
rect 2270 685 2280 735
rect 2210 675 2280 685
rect 3710 680 3730 750
rect 3800 680 4120 750
rect 3710 655 4120 680
rect 4000 588 4120 655
rect 4000 441 4121 588
rect 4000 -1509 4120 441
rect 3998 -1825 4121 -1509
rect 4000 -3291 4120 -1825
rect 3997 -3607 4121 -3291
rect 4000 -3782 4120 -3607
rect 3822 -3794 4120 -3782
rect 3822 -3894 3844 -3794
rect 3944 -3894 4120 -3794
rect 3822 -3902 4120 -3894
rect 3834 -3904 3960 -3902
<< via2 >>
rect 675 690 725 740
rect 2220 685 2270 735
rect 3844 -3894 3944 -3794
<< metal3 >>
rect 665 740 735 750
rect 665 690 675 740
rect 725 690 735 740
rect 665 680 735 690
rect 2195 735 2295 760
rect 2195 685 2220 735
rect 2270 685 2295 735
rect 2195 210 2295 685
rect 2195 110 2553 210
rect 2657 110 3828 210
rect 3728 -1920 3828 110
rect 3453 -1930 3828 -1920
rect 3453 -2030 3463 -1930
rect 3563 -2030 3828 -1930
rect 3453 -2040 3828 -2030
rect 3834 -3794 3954 -3784
rect 3834 -3894 3844 -3794
rect 3944 -3894 3954 -3794
rect 3834 -3904 3954 -3894
<< via3 >>
rect 675 690 725 740
rect 3463 -2030 3563 -1930
rect 3844 -3894 3944 -3794
<< metal4 >>
rect 665 740 735 750
rect 665 690 675 740
rect 725 690 735 740
rect 665 680 735 690
rect 675 183 725 680
rect 675 -127 725 126
rect 673 -296 726 -127
rect 3453 -1930 3573 -1920
rect 3453 -2030 3463 -1930
rect 3563 -2030 3573 -1930
rect 3453 -2040 3573 -2030
rect 3834 -3794 3954 -3784
rect 3743 -3798 3844 -3794
rect 3560 -3900 3661 -3798
rect 3693 -3894 3844 -3798
rect 3944 -3894 3954 -3794
rect 3693 -3900 3954 -3894
rect 3743 -3901 3954 -3900
rect 3822 -3904 3954 -3901
rect 3822 -3907 3944 -3904
use ro_var_extend  ro_var_extend_0
timestamp 1640959680
transform 1 0 487 0 1 675
box -375 -595 3780 765
use cbank_smol  cbank_0
timestamp 1712761727
transform 1 0 -42 0 1 -935
box 686 -840 3611 695
use cbank_smol  cbank_2
timestamp 1712761727
transform 1 0 -42 0 1 -4490
box 686 -840 3611 695
use cbank_smol  cbank_1
timestamp 1712761727
transform 1 0 -42 0 1 -2705
box 686 -840 3611 695
<< labels >>
rlabel locali 1123 -825 1123 -825 1 a0
rlabel locali 1617 -830 1617 -830 1 a1
rlabel locali 3673 -825 3673 -825 1 a5
rlabel locali 3072 -825 3072 -825 1 a4
rlabel locali 2591 -825 2591 -825 1 a3
rlabel locali 2101 -835 2101 -835 1 a2
rlabel locali 3630 370 3630 370 1 vcont
rlabel space 1275 1115 1275 1115 1 vdd!
rlabel locali 3644 713 3644 713 1 out
<< end >>
